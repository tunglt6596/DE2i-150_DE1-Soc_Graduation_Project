-- gaussian_ip_GN.vhd

-- Generated using ACDS version 17.1 590

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity gaussian_ip_GN is
	port (
		sink_data1   : in  std_logic_vector(7 downto 0) := (others => '0'); --   sink_data1.wire
		sink_eop1    : in  std_logic                    := '0';             --    sink_eop1.wire
		sink_eop2    : in  std_logic                    := '0';             --    sink_eop2.wire
		sink_valid1  : in  std_logic                    := '0';             --  sink_valid1.wire
		source_valid : out std_logic;                                       -- source_valid.wire
		sink_ready1  : out std_logic;                                       --  sink_ready1.wire
		sink_sop1    : in  std_logic                    := '0';             --    sink_sop1.wire
		source_sop   : out std_logic;                                       --   source_sop.wire
		Clock        : in  std_logic                    := '0';             --        Clock.clk
		reset        : in  std_logic                    := '0';             --             .reset
		sink_data2   : in  std_logic_vector(7 downto 0) := (others => '0'); --   sink_data2.wire
		sink_sop2    : in  std_logic                    := '0';             --    sink_sop2.wire
		source_eop   : out std_logic;                                       --   source_eop.wire
		sink_ready2  : out std_logic;                                       --  sink_ready2.wire
		source_data  : out std_logic_vector(7 downto 0);                    --  source_data.wire
		source_ready : in  std_logic                    := '0';             -- source_ready.wire
		sink_valid2  : in  std_logic                    := '0'              --  sink_valid2.wire
	);
end entity gaussian_ip_GN;

architecture rtl of gaussian_ip_GN is
	component alt_dspbuilder_clock_GNN7TLRCSZ is
		port (
			aclr      : in  std_logic := 'X'; -- reset
			aclr_n    : in  std_logic := 'X'; -- reset_n
			aclr_out  : out std_logic;        -- reset
			clock     : in  std_logic := 'X'; -- clk
			clock_out : out std_logic         -- clk
		);
	end component alt_dspbuilder_clock_GNN7TLRCSZ;

	component alt_dspbuilder_port_GN37ALZBS4 is
		port (
			input  : in  std_logic := 'X'; -- wire
			output : out std_logic         -- wire
		);
	end component alt_dspbuilder_port_GN37ALZBS4;

	component alt_dspbuilder_port_GNA5S4SQDN is
		port (
			input  : in  std_logic_vector(7 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(7 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNA5S4SQDN;

	component gaussian_ip_GN_gaussian_ip_Fusion is
		port (
			Clock     : in  std_logic                    := 'X';             -- clk
			reset     : in  std_logic                    := 'X';             -- reset
			sof_out   : out std_logic_vector(0 downto 0);                    -- wire
			valid_out : out std_logic_vector(0 downto 0);                    -- wire
			pixel2_in : in  std_logic_vector(7 downto 0) := (others => 'X'); -- wire
			pixel1_in : in  std_logic_vector(7 downto 0) := (others => 'X'); -- wire
			pixel_out : out std_logic_vector(9 downto 0);                    -- wire
			eof_out   : out std_logic_vector(0 downto 0);                    -- wire
			ready2_in : out std_logic;                                       -- wire
			valid1_in : in  std_logic                    := 'X';             -- wire
			sof1_in   : in  std_logic                    := 'X';             -- wire
			eof1_in   : in  std_logic                    := 'X'              -- wire
		);
	end component gaussian_ip_GN_gaussian_ip_Fusion;

	component alt_dspbuilder_vcc_GN is
		port (
			output : out std_logic   -- wire
		);
	end component alt_dspbuilder_vcc_GN;

	component alt_dspbuilder_cast_GN5TYUPWUA is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(9 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(7 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GN5TYUPWUA;

	component alt_dspbuilder_cast_GNSB3OXIQS is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(0 downto 0) := (others => 'X'); -- wire
			output : out std_logic                                        -- wire
		);
	end component alt_dspbuilder_cast_GNSB3OXIQS;

	signal sink_data1_0_output_wire            : std_logic_vector(7 downto 0); -- sink_data1_0:output -> gaussian_ip_Fusion_0:pixel1_in
	signal sink_data2_0_output_wire            : std_logic_vector(7 downto 0); -- sink_data2_0:output -> gaussian_ip_Fusion_0:pixel2_in
	signal sink_eop1_0_output_wire             : std_logic;                    -- sink_eop1_0:output -> gaussian_ip_Fusion_0:eof1_in
	signal vcc_output_wire                     : std_logic;                    -- VCC:output -> sink_ready1_0:input
	signal gaussian_ip_fusion_0_ready2_in_wire : std_logic;                    -- gaussian_ip_Fusion_0:ready2_in -> sink_ready2_0:input
	signal sink_sop1_0_output_wire             : std_logic;                    -- sink_sop1_0:output -> gaussian_ip_Fusion_0:sof1_in
	signal sink_valid1_0_output_wire           : std_logic;                    -- sink_valid1_0:output -> gaussian_ip_Fusion_0:valid1_in
	signal gaussian_ip_fusion_0_pixel_out_wire : std_logic_vector(9 downto 0); -- gaussian_ip_Fusion_0:pixel_out -> cast174:input
	signal cast174_output_wire                 : std_logic_vector(7 downto 0); -- cast174:output -> source_data_0:input
	signal gaussian_ip_fusion_0_eof_out_wire   : std_logic_vector(0 downto 0); -- gaussian_ip_Fusion_0:eof_out -> cast175:input
	signal cast175_output_wire                 : std_logic;                    -- cast175:output -> source_eop_0:input
	signal gaussian_ip_fusion_0_sof_out_wire   : std_logic_vector(0 downto 0); -- gaussian_ip_Fusion_0:sof_out -> cast176:input
	signal cast176_output_wire                 : std_logic;                    -- cast176:output -> source_sop_0:input
	signal gaussian_ip_fusion_0_valid_out_wire : std_logic_vector(0 downto 0); -- gaussian_ip_Fusion_0:valid_out -> cast177:input
	signal cast177_output_wire                 : std_logic;                    -- cast177:output -> source_valid_0:input
	signal clock_0_clock_output_clk            : std_logic;                    -- Clock_0:clock_out -> gaussian_ip_Fusion_0:Clock
	signal clock_0_clock_output_reset          : std_logic;                    -- Clock_0:aclr_out -> gaussian_ip_Fusion_0:reset

begin

	clock_0 : component alt_dspbuilder_clock_GNN7TLRCSZ
		port map (
			clock_out => clock_0_clock_output_clk,   -- clock_output.clk
			aclr_out  => clock_0_clock_output_reset, --             .reset
			clock     => Clock,                      --        clock.clk
			aclr      => reset                       --             .reset
		);

	source_ready_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => source_ready, --  input.wire
			output => open          -- output.wire
		);

	sink_sop1_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => sink_sop1,               --  input.wire
			output => sink_sop1_0_output_wire  -- output.wire
		);

	sink_sop2_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => sink_sop2, --  input.wire
			output => open       -- output.wire
		);

	sink_data2_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => sink_data2,               --  input.wire
			output => sink_data2_0_output_wire  -- output.wire
		);

	sink_ready1_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => vcc_output_wire, --  input.wire
			output => sink_ready1      -- output.wire
		);

	sink_data1_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => sink_data1,               --  input.wire
			output => sink_data1_0_output_wire  -- output.wire
		);

	sink_ready2_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => gaussian_ip_fusion_0_ready2_in_wire, --  input.wire
			output => sink_ready2                          -- output.wire
		);

	sink_eop1_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => sink_eop1,               --  input.wire
			output => sink_eop1_0_output_wire  -- output.wire
		);

	sink_valid2_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => sink_valid2, --  input.wire
			output => open         -- output.wire
		);

	sink_valid1_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => sink_valid1,               --  input.wire
			output => sink_valid1_0_output_wire  -- output.wire
		);

	sink_eop2_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => sink_eop2, --  input.wire
			output => open       -- output.wire
		);

	source_data_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => cast174_output_wire, --  input.wire
			output => source_data          -- output.wire
		);

	gaussian_ip_fusion_0 : component gaussian_ip_GN_gaussian_ip_Fusion
		port map (
			Clock     => clock_0_clock_output_clk,            --     Clock.clk
			reset     => clock_0_clock_output_reset,          --          .reset
			sof_out   => gaussian_ip_fusion_0_sof_out_wire,   --   sof_out.wire
			valid_out => gaussian_ip_fusion_0_valid_out_wire, -- valid_out.wire
			pixel2_in => sink_data2_0_output_wire,            -- pixel2_in.wire
			pixel1_in => sink_data1_0_output_wire,            -- pixel1_in.wire
			pixel_out => gaussian_ip_fusion_0_pixel_out_wire, -- pixel_out.wire
			eof_out   => gaussian_ip_fusion_0_eof_out_wire,   --   eof_out.wire
			ready2_in => gaussian_ip_fusion_0_ready2_in_wire, -- ready2_in.wire
			valid1_in => sink_valid1_0_output_wire,           -- valid1_in.wire
			sof1_in   => sink_sop1_0_output_wire,             --   sof1_in.wire
			eof1_in   => sink_eop1_0_output_wire              --   eof1_in.wire
		);

	source_eop_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => cast175_output_wire, --  input.wire
			output => source_eop           -- output.wire
		);

	source_valid_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => cast177_output_wire, --  input.wire
			output => source_valid         -- output.wire
		);

	source_sop_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => cast176_output_wire, --  input.wire
			output => source_sop           -- output.wire
		);

	vcc : component alt_dspbuilder_vcc_GN
		port map (
			output => vcc_output_wire  -- output.wire
		);

	cast174 : component alt_dspbuilder_cast_GN5TYUPWUA
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => gaussian_ip_fusion_0_pixel_out_wire, --  input.wire
			output => cast174_output_wire                  -- output.wire
		);

	cast175 : component alt_dspbuilder_cast_GNSB3OXIQS
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => gaussian_ip_fusion_0_eof_out_wire, --  input.wire
			output => cast175_output_wire                -- output.wire
		);

	cast176 : component alt_dspbuilder_cast_GNSB3OXIQS
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => gaussian_ip_fusion_0_sof_out_wire, --  input.wire
			output => cast176_output_wire                -- output.wire
		);

	cast177 : component alt_dspbuilder_cast_GNSB3OXIQS
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => gaussian_ip_fusion_0_valid_out_wire, --  input.wire
			output => cast177_output_wire                  -- output.wire
		);

end architecture rtl; -- of gaussian_ip_GN
