-- localedgepreserve_GN_localedgepreserve_Fusion_Cal_A_B_1_Cal_MeanI_VarI.vhd

-- Generated using ACDS version 17.1 590

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity localedgepreserve_GN_localedgepreserve_Fusion_Cal_A_B_1_Cal_MeanI_VarI is
	port (
		valid_in  : in  std_logic                     := '0';             --  valid_in.wire
		varI      : out std_logic_vector(39 downto 0);                    --      varI.wire
		Clock     : in  std_logic                     := '0';             --     Clock.clk
		reset     : in  std_logic                     := '0';             --          .reset
		pixel_in  : in  std_logic_vector(7 downto 0)  := (others => '0'); --  pixel_in.wire
		pixel_out : out std_logic_vector(7 downto 0);                     -- pixel_out.wire
		meanI     : out std_logic_vector(31 downto 0)                     --     meanI.wire
	);
end entity localedgepreserve_GN_localedgepreserve_Fusion_Cal_A_B_1_Cal_MeanI_VarI;

architecture rtl of localedgepreserve_GN_localedgepreserve_Fusion_Cal_A_B_1_Cal_MeanI_VarI is
	component alt_dspbuilder_clock_GNQFU4PUDH is
		port (
			aclr      : in  std_logic := 'X'; -- reset
			aclr_n    : in  std_logic := 'X'; -- reset_n
			aclr_out  : out std_logic;        -- reset
			clock     : in  std_logic := 'X'; -- clk
			clock_out : out std_logic         -- clk
		);
	end component alt_dspbuilder_clock_GNQFU4PUDH;

	component alt_dspbuilder_multiplier_GN64HZKYCA is
		generic (
			aWidth                         : natural := 8;
			Signed                         : natural := 0;
			bWidth                         : natural := 8;
			DEDICATED_MULTIPLIER_CIRCUITRY : string  := "AUTO";
			pipeline                       : integer := 0;
			OutputLsb                      : integer := 0;
			OutputMsb                      : integer := 8
		);
		port (
			aclr      : in  std_logic                                          := 'X';             -- clk
			clock     : in  std_logic                                          := 'X';             -- clk
			dataa     : in  std_logic_vector(aWidth-1 downto 0)                := (others => 'X'); -- wire
			datab     : in  std_logic_vector(bWidth-1 downto 0)                := (others => 'X'); -- wire
			ena       : in  std_logic                                          := 'X';             -- wire
			result    : out std_logic_vector(OutputMsb-OutputLsb+1-1 downto 0);                    -- wire
			user_aclr : in  std_logic                                          := 'X'              -- wire
		);
	end component alt_dspbuilder_multiplier_GN64HZKYCA;

	component alt_dspbuilder_gnd_GN is
		port (
			output : out std_logic   -- wire
		);
	end component alt_dspbuilder_gnd_GN;

	component alt_dspbuilder_port_GN37ALZBS4 is
		port (
			input  : in  std_logic := 'X'; -- wire
			output : out std_logic         -- wire
		);
	end component alt_dspbuilder_port_GN37ALZBS4;

	component alt_dspbuilder_multiplier_GNWZAKUPA4 is
		generic (
			aWidth                         : natural := 8;
			Signed                         : natural := 0;
			bWidth                         : natural := 8;
			DEDICATED_MULTIPLIER_CIRCUITRY : string  := "AUTO";
			pipeline                       : integer := 0;
			OutputLsb                      : integer := 0;
			OutputMsb                      : integer := 8
		);
		port (
			aclr      : in  std_logic                                          := 'X';             -- clk
			clock     : in  std_logic                                          := 'X';             -- clk
			dataa     : in  std_logic_vector(aWidth-1 downto 0)                := (others => 'X'); -- wire
			datab     : in  std_logic_vector(bWidth-1 downto 0)                := (others => 'X'); -- wire
			ena       : in  std_logic                                          := 'X';             -- wire
			result    : out std_logic_vector(OutputMsb-OutputLsb+1-1 downto 0);                    -- wire
			user_aclr : in  std_logic                                          := 'X'              -- wire
		);
	end component alt_dspbuilder_multiplier_GNWZAKUPA4;

	component alt_dspbuilder_port_GNU6ZT2WRZ is
		port (
			input  : in  std_logic_vector(39 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(39 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNU6ZT2WRZ;

	component alt_dspbuilder_memdelay_GNXMJOJMJV is
		generic (
			RAMTYPE : string   := "AUTO";
			WIDTH   : positive := 8;
			DELAY   : positive := 1
		);
		port (
			aclr      : in  std_logic                          := 'X';             -- clk
			clock     : in  std_logic                          := 'X';             -- clk
			ena       : in  std_logic                          := 'X';             -- wire
			input     : in  std_logic_vector(WIDTH-1 downto 0) := (others => 'X'); -- wire
			output    : out std_logic_vector(WIDTH-1 downto 0);                    -- wire
			user_aclr : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_memdelay_GNXMJOJMJV;

	component alt_dspbuilder_port_GNA5S4SQDN is
		port (
			input  : in  std_logic_vector(7 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(7 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNA5S4SQDN;

	component localedgepreserve_GN_localedgepreserve_Fusion_Cal_A_B_1_Cal_MeanI_VarI_MeanI is
		port (
			pixel_out : out std_logic_vector(7 downto 0);                     -- wire
			mean      : out std_logic_vector(31 downto 0);                    -- wire
			Clock     : in  std_logic                     := 'X';             -- clk
			reset     : in  std_logic                     := 'X';             -- reset
			valid_in  : in  std_logic                     := 'X';             -- wire
			pixel_in  : in  std_logic_vector(7 downto 0)  := (others => 'X')  -- wire
		);
	end component localedgepreserve_GN_localedgepreserve_Fusion_Cal_A_B_1_Cal_MeanI_VarI_MeanI;

	component alt_dspbuilder_pipelined_adder_GNY2JEH574 is
		generic (
			pipeline : integer := 0;
			width    : natural := 0
		);
		port (
			aclr      : in  std_logic                          := 'X';             -- clk
			add_sub   : in  std_logic                          := 'X';             -- wire
			cin       : in  std_logic                          := 'X';             -- wire
			clock     : in  std_logic                          := 'X';             -- clk
			cout      : out std_logic;                                             -- wire
			dataa     : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			datab     : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			ena       : in  std_logic                          := 'X';             -- wire
			result    : out std_logic_vector(width-1 downto 0);                    -- wire
			user_aclr : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_pipelined_adder_GNY2JEH574;

	component alt_dspbuilder_memdelay_GNC4CQZXMX is
		generic (
			RAMTYPE : string   := "AUTO";
			WIDTH   : positive := 8;
			DELAY   : positive := 1
		);
		port (
			aclr      : in  std_logic                          := 'X';             -- clk
			clock     : in  std_logic                          := 'X';             -- clk
			ena       : in  std_logic                          := 'X';             -- wire
			input     : in  std_logic_vector(WIDTH-1 downto 0) := (others => 'X'); -- wire
			output    : out std_logic_vector(WIDTH-1 downto 0);                    -- wire
			user_aclr : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_memdelay_GNC4CQZXMX;

	component localedgepreserve_GN_localedgepreserve_Fusion_Cal_A_B_1_Cal_MeanI_VarI_CorrI is
		port (
			corr     : out std_logic_vector(39 downto 0);                    -- wire
			Clock    : in  std_logic                     := 'X';             -- clk
			reset    : in  std_logic                     := 'X';             -- reset
			valid_in : in  std_logic                     := 'X';             -- wire
			pixel_in : in  std_logic_vector(15 downto 0) := (others => 'X')  -- wire
		);
	end component localedgepreserve_GN_localedgepreserve_Fusion_Cal_A_B_1_Cal_MeanI_VarI_CorrI;

	component alt_dspbuilder_port_GNEPKLLZKY is
		port (
			input  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(31 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNEPKLLZKY;

	component alt_dspbuilder_cast_GNR4R6OFXK is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(39 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(39 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNR4R6OFXK;

	signal multiplier2user_aclrgnd_output_wire                                      : std_logic;                     -- Multiplier2user_aclrGND:output -> Multiplier2:user_aclr
	signal multiplier1user_aclrgnd_output_wire                                      : std_logic;                     -- Multiplier1user_aclrGND:output -> Multiplier1:user_aclr
	signal memory_delay1user_aclrgnd_output_wire                                    : std_logic;                     -- Memory_Delay1user_aclrGND:output -> Memory_Delay1:user_aclr
	signal pipelined_adderuser_aclrgnd_output_wire                                  : std_logic;                     -- Pipelined_Adderuser_aclrGND:output -> Pipelined_Adder:user_aclr
	signal memory_delayuser_aclrgnd_output_wire                                     : std_logic;                     -- Memory_Delayuser_aclrGND:output -> Memory_Delay:user_aclr
	signal valid_in_0_output_wire                                                   : std_logic;                     -- valid_in_0:output -> [Memory_Delay1:ena, Memory_Delay:ena, Multiplier1:ena, Multiplier2:ena, Pipelined_Adder:ena, localedgepreserve_Fusion_Cal_A_B_1_Cal_MeanI_VarI_CorrI_0:valid_in, localedgepreserve_Fusion_Cal_A_B_1_Cal_MeanI_VarI_MeanI_0:valid_in]
	signal pixel_in_0_output_wire                                                   : std_logic_vector(7 downto 0);  -- pixel_in_0:output -> [Multiplier2:dataa, Multiplier2:datab, localedgepreserve_Fusion_Cal_A_B_1_Cal_MeanI_VarI_MeanI_0:pixel_in]
	signal localedgepreserve_fusion_cal_a_b_1_cal_meani_vari_meani_0_mean_wire      : std_logic_vector(31 downto 0); -- localedgepreserve_Fusion_Cal_A_B_1_Cal_MeanI_VarI_MeanI_0:mean -> [Memory_Delay:input, Multiplier1:dataa, Multiplier1:datab]
	signal localedgepreserve_fusion_cal_a_b_1_cal_meani_vari_meani_0_pixel_out_wire : std_logic_vector(7 downto 0);  -- localedgepreserve_Fusion_Cal_A_B_1_Cal_MeanI_VarI_MeanI_0:pixel_out -> Memory_Delay1:input
	signal multiplier2_result_wire                                                  : std_logic_vector(15 downto 0); -- Multiplier2:result -> localedgepreserve_Fusion_Cal_A_B_1_Cal_MeanI_VarI_CorrI_0:pixel_in
	signal memory_delay1_output_wire                                                : std_logic_vector(7 downto 0);  -- Memory_Delay1:output -> pixel_out_0:input
	signal pipelined_adder_result_wire                                              : std_logic_vector(39 downto 0); -- Pipelined_Adder:result -> varI_0:input
	signal memory_delay_output_wire                                                 : std_logic_vector(31 downto 0); -- Memory_Delay:output -> meanI_0:input
	signal localedgepreserve_fusion_cal_a_b_1_cal_meani_vari_corri_0_corr_wire      : std_logic_vector(39 downto 0); -- localedgepreserve_Fusion_Cal_A_B_1_Cal_MeanI_VarI_CorrI_0:corr -> cast148:input
	signal cast148_output_wire                                                      : std_logic_vector(39 downto 0); -- cast148:output -> Pipelined_Adder:dataa
	signal multiplier1_result_wire                                                  : std_logic_vector(39 downto 0); -- Multiplier1:result -> cast149:input
	signal cast149_output_wire                                                      : std_logic_vector(39 downto 0); -- cast149:output -> Pipelined_Adder:datab
	signal clock_0_clock_output_clk                                                 : std_logic;                     -- Clock_0:clock_out -> [Memory_Delay1:clock, Memory_Delay:clock, Multiplier1:clock, Multiplier2:clock, Pipelined_Adder:clock, localedgepreserve_Fusion_Cal_A_B_1_Cal_MeanI_VarI_CorrI_0:Clock, localedgepreserve_Fusion_Cal_A_B_1_Cal_MeanI_VarI_MeanI_0:Clock]
	signal clock_0_clock_output_reset                                               : std_logic;                     -- Clock_0:aclr_out -> [Memory_Delay1:aclr, Memory_Delay:aclr, Multiplier1:aclr, Multiplier2:aclr, Pipelined_Adder:aclr, localedgepreserve_Fusion_Cal_A_B_1_Cal_MeanI_VarI_CorrI_0:reset, localedgepreserve_Fusion_Cal_A_B_1_Cal_MeanI_VarI_MeanI_0:reset]

begin

	clock_0 : component alt_dspbuilder_clock_GNQFU4PUDH
		port map (
			clock_out => clock_0_clock_output_clk,   -- clock_output.clk
			aclr_out  => clock_0_clock_output_reset, --             .reset
			clock     => Clock,                      --        clock.clk
			aclr      => reset                       --             .reset
		);

	multiplier2 : component alt_dspbuilder_multiplier_GN64HZKYCA
		generic map (
			aWidth                         => 8,
			Signed                         => 0,
			bWidth                         => 8,
			DEDICATED_MULTIPLIER_CIRCUITRY => "YES",
			pipeline                       => 1,
			OutputLsb                      => 0,
			OutputMsb                      => 15
		)
		port map (
			clock     => clock_0_clock_output_clk,            -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,          --           .reset
			dataa     => pixel_in_0_output_wire,              --      dataa.wire
			datab     => pixel_in_0_output_wire,              --      datab.wire
			result    => multiplier2_result_wire,             --     result.wire
			user_aclr => multiplier2user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => valid_in_0_output_wire               --        ena.wire
		);

	multiplier2user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplier2user_aclrgnd_output_wire  -- output.wire
		);

	valid_in_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => valid_in,               --  input.wire
			output => valid_in_0_output_wire  -- output.wire
		);

	multiplier1 : component alt_dspbuilder_multiplier_GNWZAKUPA4
		generic map (
			aWidth                         => 32,
			Signed                         => 0,
			bWidth                         => 32,
			DEDICATED_MULTIPLIER_CIRCUITRY => "YES",
			pipeline                       => 1,
			OutputLsb                      => 24,
			OutputMsb                      => 63
		)
		port map (
			clock     => clock_0_clock_output_clk,                                            -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,                                          --           .reset
			dataa     => localedgepreserve_fusion_cal_a_b_1_cal_meani_vari_meani_0_mean_wire, --      dataa.wire
			datab     => localedgepreserve_fusion_cal_a_b_1_cal_meani_vari_meani_0_mean_wire, --      datab.wire
			result    => multiplier1_result_wire,                                             --     result.wire
			user_aclr => multiplier1user_aclrgnd_output_wire,                                 --  user_aclr.wire
			ena       => valid_in_0_output_wire                                               --        ena.wire
		);

	multiplier1user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplier1user_aclrgnd_output_wire  -- output.wire
		);

	vari_0 : component alt_dspbuilder_port_GNU6ZT2WRZ
		port map (
			input  => pipelined_adder_result_wire, --  input.wire
			output => varI                         -- output.wire
		);

	memory_delay1 : component alt_dspbuilder_memdelay_GNXMJOJMJV
		generic map (
			RAMTYPE => "AUTO",
			WIDTH   => 8,
			DELAY   => 2
		)
		port map (
			clock     => clock_0_clock_output_clk,                                                 -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,                                               --           .reset
			input     => localedgepreserve_fusion_cal_a_b_1_cal_meani_vari_meani_0_pixel_out_wire, --      input.wire
			output    => memory_delay1_output_wire,                                                --     output.wire
			user_aclr => memory_delay1user_aclrgnd_output_wire,                                    --  user_aclr.wire
			ena       => valid_in_0_output_wire                                                    --        ena.wire
		);

	memory_delay1user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => memory_delay1user_aclrgnd_output_wire  -- output.wire
		);

	pixel_in_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => pixel_in,               --  input.wire
			output => pixel_in_0_output_wire  -- output.wire
		);

	localedgepreserve_fusion_cal_a_b_1_cal_meani_vari_meani_0 : component localedgepreserve_GN_localedgepreserve_Fusion_Cal_A_B_1_Cal_MeanI_VarI_MeanI
		port map (
			pixel_out => localedgepreserve_fusion_cal_a_b_1_cal_meani_vari_meani_0_pixel_out_wire, -- pixel_out.wire
			mean      => localedgepreserve_fusion_cal_a_b_1_cal_meani_vari_meani_0_mean_wire,      --      mean.wire
			Clock     => clock_0_clock_output_clk,                                                 --     Clock.clk
			reset     => clock_0_clock_output_reset,                                               --          .reset
			valid_in  => valid_in_0_output_wire,                                                   --  valid_in.wire
			pixel_in  => pixel_in_0_output_wire                                                    --  pixel_in.wire
		);

	pipelined_adder : component alt_dspbuilder_pipelined_adder_GNY2JEH574
		generic map (
			pipeline => 1,
			width    => 40
		)
		port map (
			clock     => clock_0_clock_output_clk,                -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,              --           .reset
			dataa     => cast148_output_wire,                     --      dataa.wire
			datab     => cast149_output_wire,                     --      datab.wire
			result    => pipelined_adder_result_wire,             --     result.wire
			user_aclr => pipelined_adderuser_aclrgnd_output_wire, --  user_aclr.wire
			ena       => valid_in_0_output_wire                   --        ena.wire
		);

	pipelined_adderuser_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => pipelined_adderuser_aclrgnd_output_wire  -- output.wire
		);

	memory_delay : component alt_dspbuilder_memdelay_GNC4CQZXMX
		generic map (
			RAMTYPE => "AUTO",
			WIDTH   => 32,
			DELAY   => 2
		)
		port map (
			clock     => clock_0_clock_output_clk,                                            -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,                                          --           .reset
			input     => localedgepreserve_fusion_cal_a_b_1_cal_meani_vari_meani_0_mean_wire, --      input.wire
			output    => memory_delay_output_wire,                                            --     output.wire
			user_aclr => memory_delayuser_aclrgnd_output_wire,                                --  user_aclr.wire
			ena       => valid_in_0_output_wire                                               --        ena.wire
		);

	memory_delayuser_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => memory_delayuser_aclrgnd_output_wire  -- output.wire
		);

	pixel_out_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => memory_delay1_output_wire, --  input.wire
			output => pixel_out                  -- output.wire
		);

	localedgepreserve_fusion_cal_a_b_1_cal_meani_vari_corri_0 : component localedgepreserve_GN_localedgepreserve_Fusion_Cal_A_B_1_Cal_MeanI_VarI_CorrI
		port map (
			corr     => localedgepreserve_fusion_cal_a_b_1_cal_meani_vari_corri_0_corr_wire, --     corr.wire
			Clock    => clock_0_clock_output_clk,                                            --    Clock.clk
			reset    => clock_0_clock_output_reset,                                          --         .reset
			valid_in => valid_in_0_output_wire,                                              -- valid_in.wire
			pixel_in => multiplier2_result_wire                                              -- pixel_in.wire
		);

	meani_0 : component alt_dspbuilder_port_GNEPKLLZKY
		port map (
			input  => memory_delay_output_wire, --  input.wire
			output => meanI                     -- output.wire
		);

	cast148 : component alt_dspbuilder_cast_GNR4R6OFXK
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => localedgepreserve_fusion_cal_a_b_1_cal_meani_vari_corri_0_corr_wire, --  input.wire
			output => cast148_output_wire                                                  -- output.wire
		);

	cast149 : component alt_dspbuilder_cast_GNR4R6OFXK
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => multiplier1_result_wire, --  input.wire
			output => cast149_output_wire      -- output.wire
		);

end architecture rtl; -- of localedgepreserve_GN_localedgepreserve_Fusion_Cal_A_B_1_Cal_MeanI_VarI
