-- gaussian_ip_GN_gaussian_ip_Fusion_Decomposition_2_multiplier_accumulator.vhd

-- Generated using ACDS version 17.1 590

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity gaussian_ip_GN_gaussian_ip_Fusion_Decomposition_2_multiplier_accumulator is
	port (
		data_30    : in  std_logic_vector(7 downto 0)  := (others => '0'); --    data_30.wire
		data_02    : in  std_logic_vector(7 downto 0)  := (others => '0'); --    data_02.wire
		data_23    : in  std_logic_vector(7 downto 0)  := (others => '0'); --    data_23.wire
		data_43    : in  std_logic_vector(7 downto 0)  := (others => '0'); --    data_43.wire
		pixel_out  : out std_logic_vector(23 downto 0);                    --  pixel_out.wire
		data_22    : in  std_logic_vector(7 downto 0)  := (others => '0'); --    data_22.wire
		data_40    : in  std_logic_vector(7 downto 0)  := (others => '0'); --    data_40.wire
		data_20    : in  std_logic_vector(7 downto 0)  := (others => '0'); --    data_20.wire
		data_42    : in  std_logic_vector(7 downto 0)  := (others => '0'); --    data_42.wire
		Clock      : in  std_logic                     := '0';             --      Clock.clk
		reset      : in  std_logic                     := '0';             --           .reset
		data_01    : in  std_logic_vector(7 downto 0)  := (others => '0'); --    data_01.wire
		data_31    : in  std_logic_vector(7 downto 0)  := (others => '0'); --    data_31.wire
		data_10    : in  std_logic_vector(7 downto 0)  := (others => '0'); --    data_10.wire
		data_13    : in  std_logic_vector(7 downto 0)  := (others => '0'); --    data_13.wire
		data_44    : in  std_logic_vector(7 downto 0)  := (others => '0'); --    data_44.wire
		pixel_diff : out std_logic_vector(9 downto 0);                     -- pixel_diff.wire
		clken      : in  std_logic                     := '0';             --      clken.wire
		data_41    : in  std_logic_vector(7 downto 0)  := (others => '0'); --    data_41.wire
		data_34    : in  std_logic_vector(7 downto 0)  := (others => '0'); --    data_34.wire
		data_04    : in  std_logic_vector(7 downto 0)  := (others => '0'); --    data_04.wire
		data_12    : in  std_logic_vector(7 downto 0)  := (others => '0'); --    data_12.wire
		data_21    : in  std_logic_vector(7 downto 0)  := (others => '0'); --    data_21.wire
		data_00    : in  std_logic_vector(7 downto 0)  := (others => '0'); --    data_00.wire
		data_14    : in  std_logic_vector(7 downto 0)  := (others => '0'); --    data_14.wire
		data_33    : in  std_logic_vector(7 downto 0)  := (others => '0'); --    data_33.wire
		data_03    : in  std_logic_vector(7 downto 0)  := (others => '0'); --    data_03.wire
		data_11    : in  std_logic_vector(7 downto 0)  := (others => '0'); --    data_11.wire
		data_24    : in  std_logic_vector(7 downto 0)  := (others => '0'); --    data_24.wire
		data_32    : in  std_logic_vector(7 downto 0)  := (others => '0')  --    data_32.wire
	);
end entity gaussian_ip_GN_gaussian_ip_Fusion_Decomposition_2_multiplier_accumulator;

architecture rtl of gaussian_ip_GN_gaussian_ip_Fusion_Decomposition_2_multiplier_accumulator is
	component alt_dspbuilder_clock_GNQFU4PUDH is
		port (
			aclr      : in  std_logic := 'X'; -- reset
			aclr_n    : in  std_logic := 'X'; -- reset_n
			aclr_out  : out std_logic;        -- reset
			clock     : in  std_logic := 'X'; -- clk
			clock_out : out std_logic         -- clk
		);
	end component alt_dspbuilder_clock_GNQFU4PUDH;

	component alt_dspbuilder_constant_GN6SFEINY6 is
		generic (
			BitPattern : string  := "0000";
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(1 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GN6SFEINY6;

	component alt_dspbuilder_constant_GNAQNCFVSG is
		generic (
			BitPattern : string  := "0000";
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(15 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GNAQNCFVSG;

	component alt_dspbuilder_delay_GNMDMEZDYK is
		generic (
			ClockPhase : string   := "1";
			BitPattern : string   := "00000001";
			width      : positive := 8;
			use_init   : natural  := 0;
			delay      : positive := 1
		);
		port (
			aclr   : in  std_logic                          := 'X';             -- clk
			clock  : in  std_logic                          := 'X';             -- clk
			ena    : in  std_logic                          := 'X';             -- wire
			input  : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(width-1 downto 0);                    -- wire
			sclr   : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_delay_GNMDMEZDYK;

	component alt_dspbuilder_gnd_GN is
		port (
			output : out std_logic   -- wire
		);
	end component alt_dspbuilder_gnd_GN;

	component alt_dspbuilder_port_GNA5S4SQDN is
		port (
			input  : in  std_logic_vector(7 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(7 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNA5S4SQDN;

	component alt_dspbuilder_logical_bus_op_GNDCD7XEX3 is
		generic (
			logical_op       : string   := "AltAND";
			lpm_width        : positive := 8;
			shift_amount     : natural  := 3;
			mask_value       : string   := "10101010";
			signextendrshift : natural  := 1
		);
		port (
			dataa  : in  std_logic_vector(lpm_width-1 downto 0) := (others => 'X'); -- wire
			result : out std_logic_vector(lpm_width-1 downto 0)                     -- wire
		);
	end component alt_dspbuilder_logical_bus_op_GNDCD7XEX3;

	component alt_dspbuilder_multiplier_GNUH534PHC is
		generic (
			aWidth                         : natural := 8;
			Signed                         : natural := 0;
			bWidth                         : natural := 8;
			DEDICATED_MULTIPLIER_CIRCUITRY : string  := "AUTO";
			pipeline                       : integer := 0;
			OutputLsb                      : integer := 0;
			OutputMsb                      : integer := 8
		);
		port (
			aclr      : in  std_logic                                          := 'X';             -- clk
			clock     : in  std_logic                                          := 'X';             -- clk
			dataa     : in  std_logic_vector(aWidth-1 downto 0)                := (others => 'X'); -- wire
			datab     : in  std_logic_vector(bWidth-1 downto 0)                := (others => 'X'); -- wire
			ena       : in  std_logic                                          := 'X';             -- wire
			result    : out std_logic_vector(OutputMsb-OutputLsb+1-1 downto 0);                    -- wire
			user_aclr : in  std_logic                                          := 'X'              -- wire
		);
	end component alt_dspbuilder_multiplier_GNUH534PHC;

	component alt_dspbuilder_bus_concat_GNKLOJ6ING is
		generic (
			widthA : natural := 8;
			widthB : natural := 8
		);
		port (
			a      : in  std_logic_vector(widthA-1 downto 0)        := (others => 'X'); -- wire
			aclr   : in  std_logic                                  := 'X';             -- clk
			b      : in  std_logic_vector(widthB-1 downto 0)        := (others => 'X'); -- wire
			clock  : in  std_logic                                  := 'X';             -- clk
			output : out std_logic_vector(widthA+widthB-1 downto 0)                     -- wire
		);
	end component alt_dspbuilder_bus_concat_GNKLOJ6ING;

	component alt_dspbuilder_logical_bus_op_GNGAQFHY4S is
		generic (
			logical_op       : string   := "AltAND";
			lpm_width        : positive := 8;
			shift_amount     : natural  := 3;
			mask_value       : string   := "10101010";
			signextendrshift : natural  := 1
		);
		port (
			dataa  : in  std_logic_vector(lpm_width-1 downto 0) := (others => 'X'); -- wire
			result : out std_logic_vector(lpm_width-1 downto 0)                     -- wire
		);
	end component alt_dspbuilder_logical_bus_op_GNGAQFHY4S;

	component alt_dspbuilder_port_GNOC3SGKQJ is
		port (
			input  : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(23 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNOC3SGKQJ;

	component alt_dspbuilder_gain_GNIIRYXGEV is
		generic (
			InputWidth : natural := 8;
			lpm        : natural := 0;
			MaskValue  : string  := "1";
			pipeline   : natural := 0;
			gain       : string  := "00000001"
		);
		port (
			clock     : in  std_logic                     := 'X';             -- clk
			aclr      : in  std_logic                     := 'X';             -- reset
			Input     : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- wire
			Output    : out std_logic_vector(12 downto 0);                    -- wire
			user_aclr : in  std_logic                     := 'X';             -- wire
			ena       : in  std_logic                     := 'X'              -- wire
		);
	end component alt_dspbuilder_gain_GNIIRYXGEV;

	component alt_dspbuilder_delay_GNSPCBEWTM is
		generic (
			ClockPhase : string   := "1";
			BitPattern : string   := "00000001";
			width      : positive := 8;
			use_init   : natural  := 0;
			delay      : positive := 1
		);
		port (
			aclr   : in  std_logic                          := 'X';             -- clk
			clock  : in  std_logic                          := 'X';             -- clk
			ena    : in  std_logic                          := 'X';             -- wire
			input  : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(width-1 downto 0);                    -- wire
			sclr   : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_delay_GNSPCBEWTM;

	component alt_dspbuilder_delay_GNHH4N4SYH is
		generic (
			ClockPhase : string   := "1";
			BitPattern : string   := "00000001";
			width      : positive := 8;
			use_init   : natural  := 0;
			delay      : positive := 1
		);
		port (
			aclr   : in  std_logic                          := 'X';             -- clk
			clock  : in  std_logic                          := 'X';             -- clk
			ena    : in  std_logic                          := 'X';             -- wire
			input  : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(width-1 downto 0);                    -- wire
			sclr   : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_delay_GNHH4N4SYH;

	component alt_dspbuilder_pipelined_adder_GNY2JEH574 is
		generic (
			pipeline : integer := 0;
			width    : natural := 0
		);
		port (
			aclr      : in  std_logic                          := 'X';             -- clk
			add_sub   : in  std_logic                          := 'X';             -- wire
			cin       : in  std_logic                          := 'X';             -- wire
			clock     : in  std_logic                          := 'X';             -- clk
			cout      : out std_logic;                                             -- wire
			dataa     : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			datab     : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			ena       : in  std_logic                          := 'X';             -- wire
			result    : out std_logic_vector(width-1 downto 0);                    -- wire
			user_aclr : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_pipelined_adder_GNY2JEH574;

	component alt_dspbuilder_port_GNSSYS4J5R is
		port (
			input  : in  std_logic_vector(9 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(9 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNSSYS4J5R;

	component alt_dspbuilder_round_GNDZO35HDL is
		generic (
			OUT_WIDTH_g     : natural := 6;
			IN_WIDTH_g      : natural := 8;
			PIPELINE_g      : natural := 0;
			ROUNDING_TYPE_g : string  := "TRUNCATE_LOW";
			SIGNED_g        : natural := 1
		);
		port (
			clk       : in  std_logic                     := 'X';             -- clk
			reset     : in  std_logic                     := 'X';             -- wire
			datain    : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			dataout   : out std_logic_vector(7 downto 0);                     -- wire
			ena       : in  std_logic                     := 'X';             -- wire
			user_aclr : in  std_logic                     := 'X'              -- wire
		);
	end component alt_dspbuilder_round_GNDZO35HDL;

	component alt_dspbuilder_vcc_GN is
		port (
			output : out std_logic   -- wire
		);
	end component alt_dspbuilder_vcc_GN;

	component alt_dspbuilder_gain_GNBM7YKIKA is
		generic (
			InputWidth : natural := 8;
			lpm        : natural := 0;
			MaskValue  : string  := "1";
			pipeline   : natural := 0;
			gain       : string  := "00000001"
		);
		port (
			clock     : in  std_logic                     := 'X';             -- clk
			aclr      : in  std_logic                     := 'X';             -- reset
			Input     : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- wire
			Output    : out std_logic_vector(14 downto 0);                    -- wire
			user_aclr : in  std_logic                     := 'X';             -- wire
			ena       : in  std_logic                     := 'X'              -- wire
		);
	end component alt_dspbuilder_gain_GNBM7YKIKA;

	component alt_dspbuilder_delay_GN2KYXQF4S is
		generic (
			ClockPhase : string   := "1";
			BitPattern : string   := "00000001";
			width      : positive := 8;
			use_init   : natural  := 0;
			delay      : positive := 1
		);
		port (
			aclr   : in  std_logic                          := 'X';             -- clk
			clock  : in  std_logic                          := 'X';             -- clk
			ena    : in  std_logic                          := 'X';             -- wire
			input  : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(width-1 downto 0);                    -- wire
			sclr   : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_delay_GN2KYXQF4S;

	component alt_dspbuilder_gain_GNVY67KVH4 is
		generic (
			InputWidth : natural := 8;
			lpm        : natural := 0;
			MaskValue  : string  := "1";
			pipeline   : natural := 0;
			gain       : string  := "00000001"
		);
		port (
			clock     : in  std_logic                     := 'X';             -- clk
			aclr      : in  std_logic                     := 'X';             -- reset
			Input     : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- wire
			Output    : out std_logic_vector(15 downto 0);                    -- wire
			user_aclr : in  std_logic                     := 'X';             -- wire
			ena       : in  std_logic                     := 'X'              -- wire
		);
	end component alt_dspbuilder_gain_GNVY67KVH4;

	component alt_dspbuilder_parallel_adder_GNRFXUS4HJ is
		generic (
			dataWidth     : positive := 8;
			direction     : string   := "+";
			MaskValue     : string   := "1";
			pipeline      : natural  := 0;
			number_inputs : positive := 2
		);
		port (
			clock     : in  std_logic                     := 'X';             -- clk
			aclr      : in  std_logic                     := 'X';             -- reset
			result    : out std_logic_vector(20 downto 0);                    -- wire
			user_aclr : in  std_logic                     := 'X';             -- wire
			ena       : in  std_logic                     := 'X';             -- wire
			data0     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- wire
			data1     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- wire
			data2     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- wire
			data3     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- wire
			data4     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- wire
			data5     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- wire
			data6     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- wire
			data7     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- wire
			data8     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- wire
			data9     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- wire
			data10    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- wire
			data11    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- wire
			data12    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- wire
			data13    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- wire
			data14    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- wire
			data15    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- wire
			data16    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- wire
			data17    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- wire
			data18    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- wire
			data19    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- wire
			data20    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- wire
			data21    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- wire
			data22    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- wire
			data23    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- wire
			data24    : in  std_logic_vector(15 downto 0) := (others => 'X')  -- wire
		);
	end component alt_dspbuilder_parallel_adder_GNRFXUS4HJ;

	component alt_dspbuilder_delay_GNALDIUCHM is
		generic (
			ClockPhase : string   := "1";
			BitPattern : string   := "00000001";
			width      : positive := 8;
			use_init   : natural  := 0;
			delay      : positive := 1
		);
		port (
			aclr   : in  std_logic                          := 'X';             -- clk
			clock  : in  std_logic                          := 'X';             -- clk
			ena    : in  std_logic                          := 'X';             -- wire
			input  : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(width-1 downto 0);                    -- wire
			sclr   : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_delay_GNALDIUCHM;

	component alt_dspbuilder_port_GN37ALZBS4 is
		port (
			input  : in  std_logic := 'X'; -- wire
			output : out std_logic         -- wire
		);
	end component alt_dspbuilder_port_GN37ALZBS4;

	component alt_dspbuilder_memdelay_GNOQUXON7R is
		generic (
			RAMTYPE : string   := "AUTO";
			WIDTH   : positive := 8;
			DELAY   : positive := 1
		);
		port (
			aclr      : in  std_logic                          := 'X';             -- clk
			clock     : in  std_logic                          := 'X';             -- clk
			ena       : in  std_logic                          := 'X';             -- wire
			input     : in  std_logic_vector(WIDTH-1 downto 0) := (others => 'X'); -- wire
			output    : out std_logic_vector(WIDTH-1 downto 0);                    -- wire
			user_aclr : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_memdelay_GNOQUXON7R;

	component alt_dspbuilder_cast_GNUW2C7J4Q is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(7 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(8 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNUW2C7J4Q;

	component alt_dspbuilder_cast_GNNDZ2WJEB is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(7 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(9 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNNDZ2WJEB;

	component alt_dspbuilder_cast_GNUJN4ENCM is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- wire
			output : out std_logic_vector(11 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNUJN4ENCM;

	component alt_dspbuilder_cast_GNBZR5PMEK is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(7 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(7 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNBZR5PMEK;

	component alt_dspbuilder_cast_GN4Q52ZVBU is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(20 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(15 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GN4Q52ZVBU;

	component alt_dspbuilder_cast_GNT75CKW5G is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- wire
			output : out std_logic_vector(15 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNT75CKW5G;

	component alt_dspbuilder_cast_GNSGOYMYTM is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- wire
			output : out std_logic_vector(15 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNSGOYMYTM;

	component alt_dspbuilder_cast_GNYETX3347 is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(12 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(15 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNYETX3347;

	component alt_dspbuilder_cast_GNPGJSMS3Z is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(11 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(15 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNPGJSMS3Z;

	component alt_dspbuilder_cast_GNZCDPTGZG is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(14 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(15 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNZCDPTGZG;

	signal delaysclrgnd_output_wire                          : std_logic;                     -- DelaysclrGND:output -> Delay:sclr
	signal multiplier24user_aclrgnd_output_wire              : std_logic;                     -- Multiplier24user_aclrGND:output -> Multiplier24:user_aclr
	signal gainuser_aclrgnd_output_wire                      : std_logic;                     -- Gainuser_aclrGND:output -> Gain:user_aclr
	signal delay20sclrgnd_output_wire                        : std_logic;                     -- Delay20sclrGND:output -> Delay20:sclr
	signal delay22sclrgnd_output_wire                        : std_logic;                     -- Delay22sclrGND:output -> Delay22:sclr
	signal delay21sclrgnd_output_wire                        : std_logic;                     -- Delay21sclrGND:output -> Delay21:sclr
	signal delay23sclrgnd_output_wire                        : std_logic;                     -- Delay23sclrGND:output -> Delay23:sclr
	signal pipelined_adderuser_aclrgnd_output_wire           : std_logic;                     -- Pipelined_Adderuser_aclrGND:output -> Pipelined_Adder:user_aclr
	signal rounduser_aclrgnd_output_wire                     : std_logic;                     -- Rounduser_aclrGND:output -> Round:user_aclr
	signal roundenavcc_output_wire                           : std_logic;                     -- RoundenaVCC:output -> Round:ena
	signal roundresetgnd_output_wire                         : std_logic;                     -- RoundresetGND:output -> Round:reset
	signal gain5user_aclrgnd_output_wire                     : std_logic;                     -- Gain5user_aclrGND:output -> Gain5:user_aclr
	signal gain6user_aclrgnd_output_wire                     : std_logic;                     -- Gain6user_aclrGND:output -> Gain6:user_aclr
	signal delay11sclrgnd_output_wire                        : std_logic;                     -- Delay11sclrGND:output -> Delay11:sclr
	signal gain3user_aclrgnd_output_wire                     : std_logic;                     -- Gain3user_aclrGND:output -> Gain3:user_aclr
	signal delay10sclrgnd_output_wire                        : std_logic;                     -- Delay10sclrGND:output -> Delay10:sclr
	signal gain4user_aclrgnd_output_wire                     : std_logic;                     -- Gain4user_aclrGND:output -> Gain4:user_aclr
	signal delay13sclrgnd_output_wire                        : std_logic;                     -- Delay13sclrGND:output -> Delay13:sclr
	signal delay2sclrgnd_output_wire                         : std_logic;                     -- Delay2sclrGND:output -> Delay2:sclr
	signal gain1user_aclrgnd_output_wire                     : std_logic;                     -- Gain1user_aclrGND:output -> Gain1:user_aclr
	signal parallel_adder_subtractoruser_aclrgnd_output_wire : std_logic;                     -- Parallel_Adder_Subtractoruser_aclrGND:output -> Parallel_Adder_Subtractor:user_aclr
	signal delay1sclrgnd_output_wire                         : std_logic;                     -- Delay1sclrGND:output -> Delay1:sclr
	signal delay12sclrgnd_output_wire                        : std_logic;                     -- Delay12sclrGND:output -> Delay12:sclr
	signal gain2user_aclrgnd_output_wire                     : std_logic;                     -- Gain2user_aclrGND:output -> Gain2:user_aclr
	signal delay15sclrgnd_output_wire                        : std_logic;                     -- Delay15sclrGND:output -> Delay15:sclr
	signal delay14sclrgnd_output_wire                        : std_logic;                     -- Delay14sclrGND:output -> Delay14:sclr
	signal delay17sclrgnd_output_wire                        : std_logic;                     -- Delay17sclrGND:output -> Delay17:sclr
	signal delay16sclrgnd_output_wire                        : std_logic;                     -- Delay16sclrGND:output -> Delay16:sclr
	signal delay19sclrgnd_output_wire                        : std_logic;                     -- Delay19sclrGND:output -> Delay19:sclr
	signal delay18sclrgnd_output_wire                        : std_logic;                     -- Delay18sclrGND:output -> Delay18:sclr
	signal gain7user_aclrgnd_output_wire                     : std_logic;                     -- Gain7user_aclrGND:output -> Gain7:user_aclr
	signal gain8user_aclrgnd_output_wire                     : std_logic;                     -- Gain8user_aclrGND:output -> Gain8:user_aclr
	signal delay6sclrgnd_output_wire                         : std_logic;                     -- Delay6sclrGND:output -> Delay6:sclr
	signal delay5sclrgnd_output_wire                         : std_logic;                     -- Delay5sclrGND:output -> Delay5:sclr
	signal memory_delayuser_aclrgnd_output_wire              : std_logic;                     -- Memory_Delayuser_aclrGND:output -> Memory_Delay:user_aclr
	signal delay4sclrgnd_output_wire                         : std_logic;                     -- Delay4sclrGND:output -> Delay4:sclr
	signal delay3sclrgnd_output_wire                         : std_logic;                     -- Delay3sclrGND:output -> Delay3:sclr
	signal delay9sclrgnd_output_wire                         : std_logic;                     -- Delay9sclrGND:output -> Delay9:sclr
	signal delay8sclrgnd_output_wire                         : std_logic;                     -- Delay8sclrGND:output -> Delay8:sclr
	signal delay7sclrgnd_output_wire                         : std_logic;                     -- Delay7sclrGND:output -> Delay7:sclr
	signal constant25_output_wire                            : std_logic_vector(1 downto 0);  -- Constant25:output -> Bus_Concatenation1:a
	signal constant26_output_wire                            : std_logic_vector(1 downto 0);  -- Constant26:output -> Bus_Concatenation:a
	signal data_00_0_output_wire                             : std_logic_vector(7 downto 0);  -- data_00_0:output -> Delay:input
	signal data_40_0_output_wire                             : std_logic_vector(7 downto 0);  -- data_40_0:output -> Delay19:input
	signal data_04_0_output_wire                             : std_logic_vector(7 downto 0);  -- data_04_0:output -> Delay4:input
	signal clken_0_output_wire                               : std_logic;                     -- clken_0:output -> [Delay10:ena, Delay11:ena, Delay12:ena, Delay13:ena, Delay14:ena, Delay15:ena, Delay16:ena, Delay17:ena, Delay18:ena, Delay19:ena, Delay1:ena, Delay20:ena, Delay21:ena, Delay22:ena, Delay23:ena, Delay2:ena, Delay3:ena, Delay4:ena, Delay5:ena, Delay6:ena, Delay7:ena, Delay8:ena, Delay9:ena, Delay:ena, Gain1:ena, Gain2:ena, Gain3:ena, Gain4:ena, Gain5:ena, Gain6:ena, Gain7:ena, Gain8:ena, Gain:ena, Memory_Delay:ena, Multiplier24:ena, Parallel_Adder_Subtractor:ena, Pipelined_Adder:ena]
	signal data_44_0_output_wire                             : std_logic_vector(7 downto 0);  -- data_44_0:output -> Delay23:input
	signal gain_output_wire                                  : std_logic_vector(12 downto 0); -- Gain:Output -> Delay2:input
	signal gain1_output_wire                                 : std_logic_vector(14 downto 0); -- Gain1:Output -> Delay7:input
	signal gain2_output_wire                                 : std_logic_vector(12 downto 0); -- Gain2:Output -> Delay10:input
	signal gain3_output_wire                                 : std_logic_vector(14 downto 0); -- Gain3:Output -> Delay11:input
	signal gain5_output_wire                                 : std_logic_vector(14 downto 0); -- Gain5:Output -> Delay13:input
	signal gain6_output_wire                                 : std_logic_vector(12 downto 0); -- Gain6:Output -> Delay14:input
	signal gain7_output_wire                                 : std_logic_vector(14 downto 0); -- Gain7:Output -> Delay16:input
	signal gain8_output_wire                                 : std_logic_vector(12 downto 0); -- Gain8:Output -> Delay21:input
	signal logical_bus_operator_result_wire                  : std_logic_vector(9 downto 0);  -- Logical_Bus_Operator:result -> Delay1:input
	signal logical_bus_operator1_result_wire                 : std_logic_vector(9 downto 0);  -- Logical_Bus_Operator1:result -> Delay3:input
	signal logical_bus_operator10_result_wire                : std_logic_vector(9 downto 0);  -- Logical_Bus_Operator10:result -> Delay20:input
	signal logical_bus_operator11_result_wire                : std_logic_vector(9 downto 0);  -- Logical_Bus_Operator11:result -> Delay22:input
	signal logical_bus_operator2_result_wire                 : std_logic_vector(9 downto 0);  -- Logical_Bus_Operator2:result -> Delay5:input
	signal logical_bus_operator3_result_wire                 : std_logic_vector(11 downto 0); -- Logical_Bus_Operator3:result -> Delay6:input
	signal logical_bus_operator4_result_wire                 : std_logic_vector(11 downto 0); -- Logical_Bus_Operator4:result -> Delay8:input
	signal logical_bus_operator5_result_wire                 : std_logic_vector(9 downto 0);  -- Logical_Bus_Operator5:result -> Delay9:input
	signal logical_bus_operator6_result_wire                 : std_logic_vector(9 downto 0);  -- Logical_Bus_Operator6:result -> Delay12:input
	signal logical_bus_operator7_result_wire                 : std_logic_vector(11 downto 0); -- Logical_Bus_Operator7:result -> Delay15:input
	signal logical_bus_operator8_result_wire                 : std_logic_vector(11 downto 0); -- Logical_Bus_Operator8:result -> Delay17:input
	signal logical_bus_operator9_result_wire                 : std_logic_vector(9 downto 0);  -- Logical_Bus_Operator9:result -> Delay18:input
	signal data_22_0_output_wire                             : std_logic_vector(7 downto 0);  -- data_22_0:output -> [Memory_Delay:input, cast137:input]
	signal constant24_output_wire                            : std_logic_vector(15 downto 0); -- Constant24:output -> Multiplier24:datab
	signal gain4_output_wire                                 : std_logic_vector(15 downto 0); -- Gain4:Output -> Parallel_Adder_Subtractor:data12
	signal bus_concatenation1_output_wire                    : std_logic_vector(9 downto 0);  -- Bus_Concatenation1:output -> Pipelined_Adder:dataa
	signal bus_concatenation_output_wire                     : std_logic_vector(9 downto 0);  -- Bus_Concatenation:output -> Pipelined_Adder:datab
	signal multiplier24_result_wire                          : std_logic_vector(23 downto 0); -- Multiplier24:result -> [Round:datain, pixel_out_0:input]
	signal pipelined_adder_result_wire                       : std_logic_vector(9 downto 0);  -- Pipelined_Adder:result -> pixel_diff_0:input
	signal data_02_0_output_wire                             : std_logic_vector(7 downto 0);  -- data_02_0:output -> cast133:input
	signal cast133_output_wire                               : std_logic_vector(8 downto 0);  -- cast133:output -> Gain:Input
	signal data_12_0_output_wire                             : std_logic_vector(7 downto 0);  -- data_12_0:output -> cast134:input
	signal cast134_output_wire                               : std_logic_vector(8 downto 0);  -- cast134:output -> Gain1:Input
	signal data_20_0_output_wire                             : std_logic_vector(7 downto 0);  -- data_20_0:output -> cast135:input
	signal cast135_output_wire                               : std_logic_vector(8 downto 0);  -- cast135:output -> Gain2:Input
	signal data_21_0_output_wire                             : std_logic_vector(7 downto 0);  -- data_21_0:output -> cast136:input
	signal cast136_output_wire                               : std_logic_vector(8 downto 0);  -- cast136:output -> Gain3:Input
	signal cast137_output_wire                               : std_logic_vector(8 downto 0);  -- cast137:output -> Gain4:Input
	signal data_23_0_output_wire                             : std_logic_vector(7 downto 0);  -- data_23_0:output -> cast138:input
	signal cast138_output_wire                               : std_logic_vector(8 downto 0);  -- cast138:output -> Gain5:Input
	signal data_24_0_output_wire                             : std_logic_vector(7 downto 0);  -- data_24_0:output -> cast139:input
	signal cast139_output_wire                               : std_logic_vector(8 downto 0);  -- cast139:output -> Gain6:Input
	signal data_32_0_output_wire                             : std_logic_vector(7 downto 0);  -- data_32_0:output -> cast140:input
	signal cast140_output_wire                               : std_logic_vector(8 downto 0);  -- cast140:output -> Gain7:Input
	signal data_42_0_output_wire                             : std_logic_vector(7 downto 0);  -- data_42_0:output -> cast141:input
	signal cast141_output_wire                               : std_logic_vector(8 downto 0);  -- cast141:output -> Gain8:Input
	signal data_01_0_output_wire                             : std_logic_vector(7 downto 0);  -- data_01_0:output -> cast142:input
	signal cast142_output_wire                               : std_logic_vector(9 downto 0);  -- cast142:output -> Logical_Bus_Operator:dataa
	signal data_03_0_output_wire                             : std_logic_vector(7 downto 0);  -- data_03_0:output -> cast143:input
	signal cast143_output_wire                               : std_logic_vector(9 downto 0);  -- cast143:output -> Logical_Bus_Operator1:dataa
	signal data_41_0_output_wire                             : std_logic_vector(7 downto 0);  -- data_41_0:output -> cast144:input
	signal cast144_output_wire                               : std_logic_vector(9 downto 0);  -- cast144:output -> Logical_Bus_Operator10:dataa
	signal data_43_0_output_wire                             : std_logic_vector(7 downto 0);  -- data_43_0:output -> cast145:input
	signal cast145_output_wire                               : std_logic_vector(9 downto 0);  -- cast145:output -> Logical_Bus_Operator11:dataa
	signal data_10_0_output_wire                             : std_logic_vector(7 downto 0);  -- data_10_0:output -> cast146:input
	signal cast146_output_wire                               : std_logic_vector(9 downto 0);  -- cast146:output -> Logical_Bus_Operator2:dataa
	signal data_11_0_output_wire                             : std_logic_vector(7 downto 0);  -- data_11_0:output -> cast147:input
	signal cast147_output_wire                               : std_logic_vector(11 downto 0); -- cast147:output -> Logical_Bus_Operator3:dataa
	signal data_13_0_output_wire                             : std_logic_vector(7 downto 0);  -- data_13_0:output -> cast148:input
	signal cast148_output_wire                               : std_logic_vector(11 downto 0); -- cast148:output -> Logical_Bus_Operator4:dataa
	signal data_14_0_output_wire                             : std_logic_vector(7 downto 0);  -- data_14_0:output -> cast149:input
	signal cast149_output_wire                               : std_logic_vector(9 downto 0);  -- cast149:output -> Logical_Bus_Operator5:dataa
	signal data_30_0_output_wire                             : std_logic_vector(7 downto 0);  -- data_30_0:output -> cast150:input
	signal cast150_output_wire                               : std_logic_vector(9 downto 0);  -- cast150:output -> Logical_Bus_Operator6:dataa
	signal data_31_0_output_wire                             : std_logic_vector(7 downto 0);  -- data_31_0:output -> cast151:input
	signal cast151_output_wire                               : std_logic_vector(11 downto 0); -- cast151:output -> Logical_Bus_Operator7:dataa
	signal data_33_0_output_wire                             : std_logic_vector(7 downto 0);  -- data_33_0:output -> cast152:input
	signal cast152_output_wire                               : std_logic_vector(11 downto 0); -- cast152:output -> Logical_Bus_Operator8:dataa
	signal data_34_0_output_wire                             : std_logic_vector(7 downto 0);  -- data_34_0:output -> cast153:input
	signal cast153_output_wire                               : std_logic_vector(9 downto 0);  -- cast153:output -> Logical_Bus_Operator9:dataa
	signal memory_delay_output_wire                          : std_logic_vector(7 downto 0);  -- Memory_Delay:output -> cast154:input
	signal cast154_output_wire                               : std_logic_vector(7 downto 0);  -- cast154:output -> Bus_Concatenation1:b
	signal parallel_adder_subtractor_result_wire             : std_logic_vector(20 downto 0); -- Parallel_Adder_Subtractor:result -> cast155:input
	signal cast155_output_wire                               : std_logic_vector(15 downto 0); -- cast155:output -> Multiplier24:dataa
	signal delay_output_wire                                 : std_logic_vector(7 downto 0);  -- Delay:output -> cast156:input
	signal cast156_output_wire                               : std_logic_vector(15 downto 0); -- cast156:output -> Parallel_Adder_Subtractor:data0
	signal delay1_output_wire                                : std_logic_vector(9 downto 0);  -- Delay1:output -> cast157:input
	signal cast157_output_wire                               : std_logic_vector(15 downto 0); -- cast157:output -> Parallel_Adder_Subtractor:data1
	signal delay2_output_wire                                : std_logic_vector(12 downto 0); -- Delay2:output -> cast158:input
	signal cast158_output_wire                               : std_logic_vector(15 downto 0); -- cast158:output -> Parallel_Adder_Subtractor:data2
	signal delay3_output_wire                                : std_logic_vector(9 downto 0);  -- Delay3:output -> cast159:input
	signal cast159_output_wire                               : std_logic_vector(15 downto 0); -- cast159:output -> Parallel_Adder_Subtractor:data3
	signal delay4_output_wire                                : std_logic_vector(7 downto 0);  -- Delay4:output -> cast160:input
	signal cast160_output_wire                               : std_logic_vector(15 downto 0); -- cast160:output -> Parallel_Adder_Subtractor:data4
	signal delay5_output_wire                                : std_logic_vector(9 downto 0);  -- Delay5:output -> cast161:input
	signal cast161_output_wire                               : std_logic_vector(15 downto 0); -- cast161:output -> Parallel_Adder_Subtractor:data5
	signal delay6_output_wire                                : std_logic_vector(11 downto 0); -- Delay6:output -> cast162:input
	signal cast162_output_wire                               : std_logic_vector(15 downto 0); -- cast162:output -> Parallel_Adder_Subtractor:data6
	signal delay7_output_wire                                : std_logic_vector(14 downto 0); -- Delay7:output -> cast163:input
	signal cast163_output_wire                               : std_logic_vector(15 downto 0); -- cast163:output -> Parallel_Adder_Subtractor:data7
	signal delay8_output_wire                                : std_logic_vector(11 downto 0); -- Delay8:output -> cast164:input
	signal cast164_output_wire                               : std_logic_vector(15 downto 0); -- cast164:output -> Parallel_Adder_Subtractor:data8
	signal delay9_output_wire                                : std_logic_vector(9 downto 0);  -- Delay9:output -> cast165:input
	signal cast165_output_wire                               : std_logic_vector(15 downto 0); -- cast165:output -> Parallel_Adder_Subtractor:data9
	signal delay10_output_wire                               : std_logic_vector(12 downto 0); -- Delay10:output -> cast166:input
	signal cast166_output_wire                               : std_logic_vector(15 downto 0); -- cast166:output -> Parallel_Adder_Subtractor:data10
	signal delay11_output_wire                               : std_logic_vector(14 downto 0); -- Delay11:output -> cast167:input
	signal cast167_output_wire                               : std_logic_vector(15 downto 0); -- cast167:output -> Parallel_Adder_Subtractor:data11
	signal delay13_output_wire                               : std_logic_vector(14 downto 0); -- Delay13:output -> cast168:input
	signal cast168_output_wire                               : std_logic_vector(15 downto 0); -- cast168:output -> Parallel_Adder_Subtractor:data13
	signal delay14_output_wire                               : std_logic_vector(12 downto 0); -- Delay14:output -> cast169:input
	signal cast169_output_wire                               : std_logic_vector(15 downto 0); -- cast169:output -> Parallel_Adder_Subtractor:data14
	signal delay12_output_wire                               : std_logic_vector(9 downto 0);  -- Delay12:output -> cast170:input
	signal cast170_output_wire                               : std_logic_vector(15 downto 0); -- cast170:output -> Parallel_Adder_Subtractor:data15
	signal delay15_output_wire                               : std_logic_vector(11 downto 0); -- Delay15:output -> cast171:input
	signal cast171_output_wire                               : std_logic_vector(15 downto 0); -- cast171:output -> Parallel_Adder_Subtractor:data16
	signal delay16_output_wire                               : std_logic_vector(14 downto 0); -- Delay16:output -> cast172:input
	signal cast172_output_wire                               : std_logic_vector(15 downto 0); -- cast172:output -> Parallel_Adder_Subtractor:data17
	signal delay17_output_wire                               : std_logic_vector(11 downto 0); -- Delay17:output -> cast173:input
	signal cast173_output_wire                               : std_logic_vector(15 downto 0); -- cast173:output -> Parallel_Adder_Subtractor:data18
	signal delay18_output_wire                               : std_logic_vector(9 downto 0);  -- Delay18:output -> cast174:input
	signal cast174_output_wire                               : std_logic_vector(15 downto 0); -- cast174:output -> Parallel_Adder_Subtractor:data19
	signal delay19_output_wire                               : std_logic_vector(7 downto 0);  -- Delay19:output -> cast175:input
	signal cast175_output_wire                               : std_logic_vector(15 downto 0); -- cast175:output -> Parallel_Adder_Subtractor:data20
	signal delay20_output_wire                               : std_logic_vector(9 downto 0);  -- Delay20:output -> cast176:input
	signal cast176_output_wire                               : std_logic_vector(15 downto 0); -- cast176:output -> Parallel_Adder_Subtractor:data21
	signal delay21_output_wire                               : std_logic_vector(12 downto 0); -- Delay21:output -> cast177:input
	signal cast177_output_wire                               : std_logic_vector(15 downto 0); -- cast177:output -> Parallel_Adder_Subtractor:data22
	signal delay22_output_wire                               : std_logic_vector(9 downto 0);  -- Delay22:output -> cast178:input
	signal cast178_output_wire                               : std_logic_vector(15 downto 0); -- cast178:output -> Parallel_Adder_Subtractor:data23
	signal delay23_output_wire                               : std_logic_vector(7 downto 0);  -- Delay23:output -> cast179:input
	signal cast179_output_wire                               : std_logic_vector(15 downto 0); -- cast179:output -> Parallel_Adder_Subtractor:data24
	signal round_dataout_wire                                : std_logic_vector(7 downto 0);  -- Round:dataout -> cast180:input
	signal cast180_output_wire                               : std_logic_vector(7 downto 0);  -- cast180:output -> Bus_Concatenation:b
	signal clock_0_clock_output_clk                          : std_logic;                     -- Clock_0:clock_out -> [Bus_Concatenation1:clock, Bus_Concatenation:clock, Delay10:clock, Delay11:clock, Delay12:clock, Delay13:clock, Delay14:clock, Delay15:clock, Delay16:clock, Delay17:clock, Delay18:clock, Delay19:clock, Delay1:clock, Delay20:clock, Delay21:clock, Delay22:clock, Delay23:clock, Delay2:clock, Delay3:clock, Delay4:clock, Delay5:clock, Delay6:clock, Delay7:clock, Delay8:clock, Delay9:clock, Delay:clock, Gain1:clock, Gain2:clock, Gain3:clock, Gain4:clock, Gain5:clock, Gain6:clock, Gain7:clock, Gain8:clock, Gain:clock, Memory_Delay:clock, Multiplier24:clock, Parallel_Adder_Subtractor:clock, Pipelined_Adder:clock, Round:clk]
	signal clock_0_clock_output_reset                        : std_logic;                     -- Clock_0:aclr_out -> [Bus_Concatenation1:aclr, Bus_Concatenation:aclr, Delay10:aclr, Delay11:aclr, Delay12:aclr, Delay13:aclr, Delay14:aclr, Delay15:aclr, Delay16:aclr, Delay17:aclr, Delay18:aclr, Delay19:aclr, Delay1:aclr, Delay20:aclr, Delay21:aclr, Delay22:aclr, Delay23:aclr, Delay2:aclr, Delay3:aclr, Delay4:aclr, Delay5:aclr, Delay6:aclr, Delay7:aclr, Delay8:aclr, Delay9:aclr, Delay:aclr, Gain1:aclr, Gain2:aclr, Gain3:aclr, Gain4:aclr, Gain5:aclr, Gain6:aclr, Gain7:aclr, Gain8:aclr, Gain:aclr, Memory_Delay:aclr, Multiplier24:aclr, Parallel_Adder_Subtractor:aclr, Pipelined_Adder:aclr, Round:reset]

begin

	clock_0 : component alt_dspbuilder_clock_GNQFU4PUDH
		port map (
			clock_out => clock_0_clock_output_clk,   -- clock_output.clk
			aclr_out  => clock_0_clock_output_reset, --             .reset
			clock     => Clock,                      --        clock.clk
			aclr      => reset                       --             .reset
		);

	constant26 : component alt_dspbuilder_constant_GN6SFEINY6
		generic map (
			BitPattern => "00",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 2
		)
		port map (
			output => constant26_output_wire  -- output.wire
		);

	constant25 : component alt_dspbuilder_constant_GN6SFEINY6
		generic map (
			BitPattern => "00",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 2
		)
		port map (
			output => constant25_output_wire  -- output.wire
		);

	constant24 : component alt_dspbuilder_constant_GNAQNCFVSG
		generic map (
			BitPattern => "0000000100000000",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 16
		)
		port map (
			output => constant24_output_wire  -- output.wire
		);

	delay : component alt_dspbuilder_delay_GNMDMEZDYK
		generic map (
			ClockPhase => "1",
			BitPattern => "00000001",
			width      => 8,
			use_init   => 0,
			delay      => 6
		)
		port map (
			input  => data_00_0_output_wire,      --      input.wire
			clock  => clock_0_clock_output_clk,   -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset, --           .reset
			output => delay_output_wire,          --     output.wire
			sclr   => delaysclrgnd_output_wire,   --       sclr.wire
			ena    => clken_0_output_wire         --        ena.wire
		);

	delaysclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delaysclrgnd_output_wire  -- output.wire
		);

	data_33_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => data_33,               --  input.wire
			output => data_33_0_output_wire  -- output.wire
		);

	data_32_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => data_32,               --  input.wire
			output => data_32_0_output_wire  -- output.wire
		);

	data_34_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => data_34,               --  input.wire
			output => data_34_0_output_wire  -- output.wire
		);

	data_31_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => data_31,               --  input.wire
			output => data_31_0_output_wire  -- output.wire
		);

	data_30_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => data_30,               --  input.wire
			output => data_30_0_output_wire  -- output.wire
		);

	logical_bus_operator : component alt_dspbuilder_logical_bus_op_GNDCD7XEX3
		generic map (
			logical_op       => "AltShiftLeft",
			lpm_width        => 10,
			shift_amount     => 2,
			mask_value       => "1111111011",
			signextendrshift => 0
		)
		port map (
			dataa  => cast142_output_wire,              --  dataa.wire
			result => logical_bus_operator_result_wire  -- result.wire
		);

	multiplier24 : component alt_dspbuilder_multiplier_GNUH534PHC
		generic map (
			aWidth                         => 16,
			Signed                         => 0,
			bWidth                         => 16,
			DEDICATED_MULTIPLIER_CIRCUITRY => "NO",
			pipeline                       => 16,
			OutputLsb                      => 0,
			OutputMsb                      => 23
		)
		port map (
			clock     => clock_0_clock_output_clk,             -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,           --           .reset
			dataa     => cast155_output_wire,                  --      dataa.wire
			datab     => constant24_output_wire,               --      datab.wire
			result    => multiplier24_result_wire,             --     result.wire
			user_aclr => multiplier24user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => clken_0_output_wire                   --        ena.wire
		);

	multiplier24user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplier24user_aclrgnd_output_wire  -- output.wire
		);

	logical_bus_operator10 : component alt_dspbuilder_logical_bus_op_GNDCD7XEX3
		generic map (
			logical_op       => "AltShiftLeft",
			lpm_width        => 10,
			shift_amount     => 2,
			mask_value       => "1111111011",
			signextendrshift => 0
		)
		port map (
			dataa  => cast144_output_wire,                --  dataa.wire
			result => logical_bus_operator10_result_wire  -- result.wire
		);

	logical_bus_operator11 : component alt_dspbuilder_logical_bus_op_GNDCD7XEX3
		generic map (
			logical_op       => "AltShiftLeft",
			lpm_width        => 10,
			shift_amount     => 2,
			mask_value       => "1111111011",
			signextendrshift => 0
		)
		port map (
			dataa  => cast145_output_wire,                --  dataa.wire
			result => logical_bus_operator11_result_wire  -- result.wire
		);

	data_00_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => data_00,               --  input.wire
			output => data_00_0_output_wire  -- output.wire
		);

	data_44_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => data_44,               --  input.wire
			output => data_44_0_output_wire  -- output.wire
		);

	bus_concatenation1 : component alt_dspbuilder_bus_concat_GNKLOJ6ING
		generic map (
			widthA => 2,
			widthB => 8
		)
		port map (
			clock  => clock_0_clock_output_clk,       -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,     --           .reset
			a      => constant25_output_wire,         --          a.wire
			b      => cast154_output_wire,            --          b.wire
			output => bus_concatenation1_output_wire  --     output.wire
		);

	logical_bus_operator8 : component alt_dspbuilder_logical_bus_op_GNGAQFHY4S
		generic map (
			logical_op       => "AltShiftLeft",
			lpm_width        => 12,
			shift_amount     => 4,
			mask_value       => "111111111011",
			signextendrshift => 0
		)
		port map (
			dataa  => cast152_output_wire,               --  dataa.wire
			result => logical_bus_operator8_result_wire  -- result.wire
		);

	data_43_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => data_43,               --  input.wire
			output => data_43_0_output_wire  -- output.wire
		);

	logical_bus_operator7 : component alt_dspbuilder_logical_bus_op_GNGAQFHY4S
		generic map (
			logical_op       => "AltShiftLeft",
			lpm_width        => 12,
			shift_amount     => 4,
			mask_value       => "111111111011",
			signextendrshift => 0
		)
		port map (
			dataa  => cast151_output_wire,               --  dataa.wire
			result => logical_bus_operator7_result_wire  -- result.wire
		);

	data_02_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => data_02,               --  input.wire
			output => data_02_0_output_wire  -- output.wire
		);

	logical_bus_operator6 : component alt_dspbuilder_logical_bus_op_GNDCD7XEX3
		generic map (
			logical_op       => "AltShiftLeft",
			lpm_width        => 10,
			shift_amount     => 2,
			mask_value       => "1111111011",
			signextendrshift => 0
		)
		port map (
			dataa  => cast150_output_wire,               --  dataa.wire
			result => logical_bus_operator6_result_wire  -- result.wire
		);

	data_01_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => data_01,               --  input.wire
			output => data_01_0_output_wire  -- output.wire
		);

	logical_bus_operator5 : component alt_dspbuilder_logical_bus_op_GNDCD7XEX3
		generic map (
			logical_op       => "AltShiftLeft",
			lpm_width        => 10,
			shift_amount     => 2,
			mask_value       => "1111111011",
			signextendrshift => 0
		)
		port map (
			dataa  => cast149_output_wire,               --  dataa.wire
			result => logical_bus_operator5_result_wire  -- result.wire
		);

	data_40_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => data_40,               --  input.wire
			output => data_40_0_output_wire  -- output.wire
		);

	logical_bus_operator4 : component alt_dspbuilder_logical_bus_op_GNGAQFHY4S
		generic map (
			logical_op       => "AltShiftLeft",
			lpm_width        => 12,
			shift_amount     => 4,
			mask_value       => "111111111011",
			signextendrshift => 0
		)
		port map (
			dataa  => cast148_output_wire,               --  dataa.wire
			result => logical_bus_operator4_result_wire  -- result.wire
		);

	logical_bus_operator3 : component alt_dspbuilder_logical_bus_op_GNGAQFHY4S
		generic map (
			logical_op       => "AltShiftLeft",
			lpm_width        => 12,
			shift_amount     => 4,
			mask_value       => "111111111011",
			signextendrshift => 0
		)
		port map (
			dataa  => cast147_output_wire,               --  dataa.wire
			result => logical_bus_operator3_result_wire  -- result.wire
		);

	data_42_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => data_42,               --  input.wire
			output => data_42_0_output_wire  -- output.wire
		);

	logical_bus_operator2 : component alt_dspbuilder_logical_bus_op_GNDCD7XEX3
		generic map (
			logical_op       => "AltShiftLeft",
			lpm_width        => 10,
			shift_amount     => 2,
			mask_value       => "1111111011",
			signextendrshift => 0
		)
		port map (
			dataa  => cast146_output_wire,               --  dataa.wire
			result => logical_bus_operator2_result_wire  -- result.wire
		);

	data_41_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => data_41,               --  input.wire
			output => data_41_0_output_wire  -- output.wire
		);

	logical_bus_operator1 : component alt_dspbuilder_logical_bus_op_GNDCD7XEX3
		generic map (
			logical_op       => "AltShiftLeft",
			lpm_width        => 10,
			shift_amount     => 2,
			mask_value       => "1111111011",
			signextendrshift => 0
		)
		port map (
			dataa  => cast143_output_wire,               --  dataa.wire
			result => logical_bus_operator1_result_wire  -- result.wire
		);

	pixel_out_0 : component alt_dspbuilder_port_GNOC3SGKQJ
		port map (
			input  => multiplier24_result_wire, --  input.wire
			output => pixel_out                 -- output.wire
		);

	data_04_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => data_04,               --  input.wire
			output => data_04_0_output_wire  -- output.wire
		);

	data_03_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => data_03,               --  input.wire
			output => data_03_0_output_wire  -- output.wire
		);

	gain : component alt_dspbuilder_gain_GNIIRYXGEV
		generic map (
			InputWidth => 9,
			lpm        => 0,
			MaskValue  => "1",
			pipeline   => 3,
			gain       => "0110"
		)
		port map (
			clock     => clock_0_clock_output_clk,     -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,   --           .reset
			Input     => cast133_output_wire,          --      Input.wire
			Output    => gain_output_wire,             --     Output.wire
			user_aclr => gainuser_aclrgnd_output_wire, --  user_aclr.wire
			ena       => clken_0_output_wire           --        ena.wire
		);

	gainuser_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => gainuser_aclrgnd_output_wire  -- output.wire
		);

	delay20 : component alt_dspbuilder_delay_GNSPCBEWTM
		generic map (
			ClockPhase => "1",
			BitPattern => "0000000001",
			width      => 10,
			use_init   => 0,
			delay      => 6
		)
		port map (
			input  => logical_bus_operator10_result_wire, --      input.wire
			clock  => clock_0_clock_output_clk,           -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,         --           .reset
			output => delay20_output_wire,                --     output.wire
			sclr   => delay20sclrgnd_output_wire,         --       sclr.wire
			ena    => clken_0_output_wire                 --        ena.wire
		);

	delay20sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delay20sclrgnd_output_wire  -- output.wire
		);

	delay22 : component alt_dspbuilder_delay_GNSPCBEWTM
		generic map (
			ClockPhase => "1",
			BitPattern => "0000000001",
			width      => 10,
			use_init   => 0,
			delay      => 6
		)
		port map (
			input  => logical_bus_operator11_result_wire, --      input.wire
			clock  => clock_0_clock_output_clk,           -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,         --           .reset
			output => delay22_output_wire,                --     output.wire
			sclr   => delay22sclrgnd_output_wire,         --       sclr.wire
			ena    => clken_0_output_wire                 --        ena.wire
		);

	delay22sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delay22sclrgnd_output_wire  -- output.wire
		);

	delay21 : component alt_dspbuilder_delay_GNHH4N4SYH
		generic map (
			ClockPhase => "1",
			BitPattern => "0000000000001",
			width      => 13,
			use_init   => 0,
			delay      => 3
		)
		port map (
			input  => gain8_output_wire,          --      input.wire
			clock  => clock_0_clock_output_clk,   -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset, --           .reset
			output => delay21_output_wire,        --     output.wire
			sclr   => delay21sclrgnd_output_wire, --       sclr.wire
			ena    => clken_0_output_wire         --        ena.wire
		);

	delay21sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delay21sclrgnd_output_wire  -- output.wire
		);

	delay23 : component alt_dspbuilder_delay_GNMDMEZDYK
		generic map (
			ClockPhase => "1",
			BitPattern => "00000001",
			width      => 8,
			use_init   => 0,
			delay      => 6
		)
		port map (
			input  => data_44_0_output_wire,      --      input.wire
			clock  => clock_0_clock_output_clk,   -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset, --           .reset
			output => delay23_output_wire,        --     output.wire
			sclr   => delay23sclrgnd_output_wire, --       sclr.wire
			ena    => clken_0_output_wire         --        ena.wire
		);

	delay23sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delay23sclrgnd_output_wire  -- output.wire
		);

	bus_concatenation : component alt_dspbuilder_bus_concat_GNKLOJ6ING
		generic map (
			widthA => 2,
			widthB => 8
		)
		port map (
			clock  => clock_0_clock_output_clk,      -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,    --           .reset
			a      => constant26_output_wire,        --          a.wire
			b      => cast180_output_wire,           --          b.wire
			output => bus_concatenation_output_wire  --     output.wire
		);

	pipelined_adder : component alt_dspbuilder_pipelined_adder_GNY2JEH574
		generic map (
			pipeline => 1,
			width    => 10
		)
		port map (
			clock     => clock_0_clock_output_clk,                -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,              --           .reset
			dataa     => bus_concatenation1_output_wire,          --      dataa.wire
			datab     => bus_concatenation_output_wire,           --      datab.wire
			result    => pipelined_adder_result_wire,             --     result.wire
			user_aclr => pipelined_adderuser_aclrgnd_output_wire, --  user_aclr.wire
			ena       => clken_0_output_wire                      --        ena.wire
		);

	pipelined_adderuser_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => pipelined_adderuser_aclrgnd_output_wire  -- output.wire
		);

	logical_bus_operator9 : component alt_dspbuilder_logical_bus_op_GNDCD7XEX3
		generic map (
			logical_op       => "AltShiftLeft",
			lpm_width        => 10,
			shift_amount     => 2,
			mask_value       => "1111111011",
			signextendrshift => 0
		)
		port map (
			dataa  => cast153_output_wire,               --  dataa.wire
			result => logical_bus_operator9_result_wire  -- result.wire
		);

	data_11_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => data_11,               --  input.wire
			output => data_11_0_output_wire  -- output.wire
		);

	data_10_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => data_10,               --  input.wire
			output => data_10_0_output_wire  -- output.wire
		);

	data_13_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => data_13,               --  input.wire
			output => data_13_0_output_wire  -- output.wire
		);

	data_12_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => data_12,               --  input.wire
			output => data_12_0_output_wire  -- output.wire
		);

	pixel_diff_0 : component alt_dspbuilder_port_GNSSYS4J5R
		port map (
			input  => pipelined_adder_result_wire, --  input.wire
			output => pixel_diff                   -- output.wire
		);

	round : component alt_dspbuilder_round_GNDZO35HDL
		generic map (
			OUT_WIDTH_g     => 8,
			IN_WIDTH_g      => 24,
			PIPELINE_g      => 0,
			ROUNDING_TYPE_g => "ROUND_UP",
			SIGNED_g        => 0
		)
		port map (
			clk       => clock_0_clock_output_clk,      -- clk_reset.clk
			reset     => clock_0_clock_output_reset,    --          .reset
			datain    => multiplier24_result_wire,      --    datain.wire
			dataout   => round_dataout_wire,            --   dataout.wire
			ena       => roundenavcc_output_wire,       --       ena.wire
			user_aclr => rounduser_aclrgnd_output_wire  -- user_aclr.wire
		);

	rounduser_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => rounduser_aclrgnd_output_wire  -- output.wire
		);

	roundenavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => roundenavcc_output_wire  -- output.wire
		);

	roundresetgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => roundresetgnd_output_wire  -- output.wire
		);

	data_14_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => data_14,               --  input.wire
			output => data_14_0_output_wire  -- output.wire
		);

	gain5 : component alt_dspbuilder_gain_GNBM7YKIKA
		generic map (
			InputWidth => 9,
			lpm        => 0,
			MaskValue  => "1",
			pipeline   => 5,
			gain       => "011000"
		)
		port map (
			clock     => clock_0_clock_output_clk,      -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,    --           .reset
			Input     => cast138_output_wire,           --      Input.wire
			Output    => gain5_output_wire,             --     Output.wire
			user_aclr => gain5user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => clken_0_output_wire            --        ena.wire
		);

	gain5user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => gain5user_aclrgnd_output_wire  -- output.wire
		);

	gain6 : component alt_dspbuilder_gain_GNIIRYXGEV
		generic map (
			InputWidth => 9,
			lpm        => 0,
			MaskValue  => "1",
			pipeline   => 3,
			gain       => "0110"
		)
		port map (
			clock     => clock_0_clock_output_clk,      -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,    --           .reset
			Input     => cast139_output_wire,           --      Input.wire
			Output    => gain6_output_wire,             --     Output.wire
			user_aclr => gain6user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => clken_0_output_wire            --        ena.wire
		);

	gain6user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => gain6user_aclrgnd_output_wire  -- output.wire
		);

	delay11 : component alt_dspbuilder_delay_GN2KYXQF4S
		generic map (
			ClockPhase => "1",
			BitPattern => "000000000000001",
			width      => 15,
			use_init   => 0,
			delay      => 1
		)
		port map (
			input  => gain3_output_wire,          --      input.wire
			clock  => clock_0_clock_output_clk,   -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset, --           .reset
			output => delay11_output_wire,        --     output.wire
			sclr   => delay11sclrgnd_output_wire, --       sclr.wire
			ena    => clken_0_output_wire         --        ena.wire
		);

	delay11sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delay11sclrgnd_output_wire  -- output.wire
		);

	gain3 : component alt_dspbuilder_gain_GNBM7YKIKA
		generic map (
			InputWidth => 9,
			lpm        => 0,
			MaskValue  => "1",
			pipeline   => 5,
			gain       => "011000"
		)
		port map (
			clock     => clock_0_clock_output_clk,      -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,    --           .reset
			Input     => cast136_output_wire,           --      Input.wire
			Output    => gain3_output_wire,             --     Output.wire
			user_aclr => gain3user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => clken_0_output_wire            --        ena.wire
		);

	gain3user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => gain3user_aclrgnd_output_wire  -- output.wire
		);

	delay10 : component alt_dspbuilder_delay_GNHH4N4SYH
		generic map (
			ClockPhase => "1",
			BitPattern => "0000000000001",
			width      => 13,
			use_init   => 0,
			delay      => 3
		)
		port map (
			input  => gain2_output_wire,          --      input.wire
			clock  => clock_0_clock_output_clk,   -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset, --           .reset
			output => delay10_output_wire,        --     output.wire
			sclr   => delay10sclrgnd_output_wire, --       sclr.wire
			ena    => clken_0_output_wire         --        ena.wire
		);

	delay10sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delay10sclrgnd_output_wire  -- output.wire
		);

	gain4 : component alt_dspbuilder_gain_GNVY67KVH4
		generic map (
			InputWidth => 9,
			lpm        => 0,
			MaskValue  => "1",
			pipeline   => 6,
			gain       => "0100100"
		)
		port map (
			clock     => clock_0_clock_output_clk,      -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,    --           .reset
			Input     => cast137_output_wire,           --      Input.wire
			Output    => gain4_output_wire,             --     Output.wire
			user_aclr => gain4user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => clken_0_output_wire            --        ena.wire
		);

	gain4user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => gain4user_aclrgnd_output_wire  -- output.wire
		);

	delay13 : component alt_dspbuilder_delay_GN2KYXQF4S
		generic map (
			ClockPhase => "1",
			BitPattern => "000000000000001",
			width      => 15,
			use_init   => 0,
			delay      => 1
		)
		port map (
			input  => gain5_output_wire,          --      input.wire
			clock  => clock_0_clock_output_clk,   -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset, --           .reset
			output => delay13_output_wire,        --     output.wire
			sclr   => delay13sclrgnd_output_wire, --       sclr.wire
			ena    => clken_0_output_wire         --        ena.wire
		);

	delay13sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delay13sclrgnd_output_wire  -- output.wire
		);

	delay2 : component alt_dspbuilder_delay_GNHH4N4SYH
		generic map (
			ClockPhase => "1",
			BitPattern => "0000000000001",
			width      => 13,
			use_init   => 0,
			delay      => 3
		)
		port map (
			input  => gain_output_wire,           --      input.wire
			clock  => clock_0_clock_output_clk,   -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset, --           .reset
			output => delay2_output_wire,         --     output.wire
			sclr   => delay2sclrgnd_output_wire,  --       sclr.wire
			ena    => clken_0_output_wire         --        ena.wire
		);

	delay2sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delay2sclrgnd_output_wire  -- output.wire
		);

	gain1 : component alt_dspbuilder_gain_GNBM7YKIKA
		generic map (
			InputWidth => 9,
			lpm        => 0,
			MaskValue  => "1",
			pipeline   => 5,
			gain       => "011000"
		)
		port map (
			clock     => clock_0_clock_output_clk,      -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,    --           .reset
			Input     => cast134_output_wire,           --      Input.wire
			Output    => gain1_output_wire,             --     Output.wire
			user_aclr => gain1user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => clken_0_output_wire            --        ena.wire
		);

	gain1user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => gain1user_aclrgnd_output_wire  -- output.wire
		);

	parallel_adder_subtractor : component alt_dspbuilder_parallel_adder_GNRFXUS4HJ
		generic map (
			dataWidth     => 16,
			direction     => "+",
			MaskValue     => "1",
			pipeline      => 1,
			number_inputs => 25
		)
		port map (
			clock     => clock_0_clock_output_clk,                          -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,                        --           .reset
			result    => parallel_adder_subtractor_result_wire,             --     result.wire
			user_aclr => parallel_adder_subtractoruser_aclrgnd_output_wire, --  user_aclr.wire
			ena       => clken_0_output_wire,                               --        ena.wire
			data0     => cast156_output_wire,                               --      data0.wire
			data1     => cast157_output_wire,                               --      data1.wire
			data2     => cast158_output_wire,                               --      data2.wire
			data3     => cast159_output_wire,                               --      data3.wire
			data4     => cast160_output_wire,                               --      data4.wire
			data5     => cast161_output_wire,                               --      data5.wire
			data6     => cast162_output_wire,                               --      data6.wire
			data7     => cast163_output_wire,                               --      data7.wire
			data8     => cast164_output_wire,                               --      data8.wire
			data9     => cast165_output_wire,                               --      data9.wire
			data10    => cast166_output_wire,                               --     data10.wire
			data11    => cast167_output_wire,                               --     data11.wire
			data12    => gain4_output_wire,                                 --     data12.wire
			data13    => cast168_output_wire,                               --     data13.wire
			data14    => cast169_output_wire,                               --     data14.wire
			data15    => cast170_output_wire,                               --     data15.wire
			data16    => cast171_output_wire,                               --     data16.wire
			data17    => cast172_output_wire,                               --     data17.wire
			data18    => cast173_output_wire,                               --     data18.wire
			data19    => cast174_output_wire,                               --     data19.wire
			data20    => cast175_output_wire,                               --     data20.wire
			data21    => cast176_output_wire,                               --     data21.wire
			data22    => cast177_output_wire,                               --     data22.wire
			data23    => cast178_output_wire,                               --     data23.wire
			data24    => cast179_output_wire                                --     data24.wire
		);

	parallel_adder_subtractoruser_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => parallel_adder_subtractoruser_aclrgnd_output_wire  -- output.wire
		);

	delay1 : component alt_dspbuilder_delay_GNSPCBEWTM
		generic map (
			ClockPhase => "1",
			BitPattern => "0000000001",
			width      => 10,
			use_init   => 0,
			delay      => 6
		)
		port map (
			input  => logical_bus_operator_result_wire, --      input.wire
			clock  => clock_0_clock_output_clk,         -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,       --           .reset
			output => delay1_output_wire,               --     output.wire
			sclr   => delay1sclrgnd_output_wire,        --       sclr.wire
			ena    => clken_0_output_wire               --        ena.wire
		);

	delay1sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delay1sclrgnd_output_wire  -- output.wire
		);

	delay12 : component alt_dspbuilder_delay_GNSPCBEWTM
		generic map (
			ClockPhase => "1",
			BitPattern => "0000000001",
			width      => 10,
			use_init   => 0,
			delay      => 6
		)
		port map (
			input  => logical_bus_operator6_result_wire, --      input.wire
			clock  => clock_0_clock_output_clk,          -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,        --           .reset
			output => delay12_output_wire,               --     output.wire
			sclr   => delay12sclrgnd_output_wire,        --       sclr.wire
			ena    => clken_0_output_wire                --        ena.wire
		);

	delay12sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delay12sclrgnd_output_wire  -- output.wire
		);

	gain2 : component alt_dspbuilder_gain_GNIIRYXGEV
		generic map (
			InputWidth => 9,
			lpm        => 0,
			MaskValue  => "1",
			pipeline   => 3,
			gain       => "0110"
		)
		port map (
			clock     => clock_0_clock_output_clk,      -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,    --           .reset
			Input     => cast135_output_wire,           --      Input.wire
			Output    => gain2_output_wire,             --     Output.wire
			user_aclr => gain2user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => clken_0_output_wire            --        ena.wire
		);

	gain2user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => gain2user_aclrgnd_output_wire  -- output.wire
		);

	delay15 : component alt_dspbuilder_delay_GNALDIUCHM
		generic map (
			ClockPhase => "1",
			BitPattern => "000000000001",
			width      => 12,
			use_init   => 0,
			delay      => 6
		)
		port map (
			input  => logical_bus_operator7_result_wire, --      input.wire
			clock  => clock_0_clock_output_clk,          -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,        --           .reset
			output => delay15_output_wire,               --     output.wire
			sclr   => delay15sclrgnd_output_wire,        --       sclr.wire
			ena    => clken_0_output_wire                --        ena.wire
		);

	delay15sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delay15sclrgnd_output_wire  -- output.wire
		);

	delay14 : component alt_dspbuilder_delay_GNHH4N4SYH
		generic map (
			ClockPhase => "1",
			BitPattern => "0000000000001",
			width      => 13,
			use_init   => 0,
			delay      => 3
		)
		port map (
			input  => gain6_output_wire,          --      input.wire
			clock  => clock_0_clock_output_clk,   -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset, --           .reset
			output => delay14_output_wire,        --     output.wire
			sclr   => delay14sclrgnd_output_wire, --       sclr.wire
			ena    => clken_0_output_wire         --        ena.wire
		);

	delay14sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delay14sclrgnd_output_wire  -- output.wire
		);

	delay17 : component alt_dspbuilder_delay_GNALDIUCHM
		generic map (
			ClockPhase => "1",
			BitPattern => "000000000001",
			width      => 12,
			use_init   => 0,
			delay      => 6
		)
		port map (
			input  => logical_bus_operator8_result_wire, --      input.wire
			clock  => clock_0_clock_output_clk,          -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,        --           .reset
			output => delay17_output_wire,               --     output.wire
			sclr   => delay17sclrgnd_output_wire,        --       sclr.wire
			ena    => clken_0_output_wire                --        ena.wire
		);

	delay17sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delay17sclrgnd_output_wire  -- output.wire
		);

	delay16 : component alt_dspbuilder_delay_GN2KYXQF4S
		generic map (
			ClockPhase => "1",
			BitPattern => "000000000000001",
			width      => 15,
			use_init   => 0,
			delay      => 1
		)
		port map (
			input  => gain7_output_wire,          --      input.wire
			clock  => clock_0_clock_output_clk,   -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset, --           .reset
			output => delay16_output_wire,        --     output.wire
			sclr   => delay16sclrgnd_output_wire, --       sclr.wire
			ena    => clken_0_output_wire         --        ena.wire
		);

	delay16sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delay16sclrgnd_output_wire  -- output.wire
		);

	delay19 : component alt_dspbuilder_delay_GNMDMEZDYK
		generic map (
			ClockPhase => "1",
			BitPattern => "00000001",
			width      => 8,
			use_init   => 0,
			delay      => 6
		)
		port map (
			input  => data_40_0_output_wire,      --      input.wire
			clock  => clock_0_clock_output_clk,   -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset, --           .reset
			output => delay19_output_wire,        --     output.wire
			sclr   => delay19sclrgnd_output_wire, --       sclr.wire
			ena    => clken_0_output_wire         --        ena.wire
		);

	delay19sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delay19sclrgnd_output_wire  -- output.wire
		);

	delay18 : component alt_dspbuilder_delay_GNSPCBEWTM
		generic map (
			ClockPhase => "1",
			BitPattern => "0000000001",
			width      => 10,
			use_init   => 0,
			delay      => 6
		)
		port map (
			input  => logical_bus_operator9_result_wire, --      input.wire
			clock  => clock_0_clock_output_clk,          -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,        --           .reset
			output => delay18_output_wire,               --     output.wire
			sclr   => delay18sclrgnd_output_wire,        --       sclr.wire
			ena    => clken_0_output_wire                --        ena.wire
		);

	delay18sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delay18sclrgnd_output_wire  -- output.wire
		);

	clken_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => clken,               --  input.wire
			output => clken_0_output_wire  -- output.wire
		);

	gain7 : component alt_dspbuilder_gain_GNBM7YKIKA
		generic map (
			InputWidth => 9,
			lpm        => 0,
			MaskValue  => "1",
			pipeline   => 5,
			gain       => "011000"
		)
		port map (
			clock     => clock_0_clock_output_clk,      -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,    --           .reset
			Input     => cast140_output_wire,           --      Input.wire
			Output    => gain7_output_wire,             --     Output.wire
			user_aclr => gain7user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => clken_0_output_wire            --        ena.wire
		);

	gain7user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => gain7user_aclrgnd_output_wire  -- output.wire
		);

	gain8 : component alt_dspbuilder_gain_GNIIRYXGEV
		generic map (
			InputWidth => 9,
			lpm        => 0,
			MaskValue  => "1",
			pipeline   => 3,
			gain       => "0110"
		)
		port map (
			clock     => clock_0_clock_output_clk,      -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,    --           .reset
			Input     => cast141_output_wire,           --      Input.wire
			Output    => gain8_output_wire,             --     Output.wire
			user_aclr => gain8user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => clken_0_output_wire            --        ena.wire
		);

	gain8user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => gain8user_aclrgnd_output_wire  -- output.wire
		);

	data_22_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => data_22,               --  input.wire
			output => data_22_0_output_wire  -- output.wire
		);

	data_21_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => data_21,               --  input.wire
			output => data_21_0_output_wire  -- output.wire
		);

	data_24_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => data_24,               --  input.wire
			output => data_24_0_output_wire  -- output.wire
		);

	data_23_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => data_23,               --  input.wire
			output => data_23_0_output_wire  -- output.wire
		);

	data_20_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => data_20,               --  input.wire
			output => data_20_0_output_wire  -- output.wire
		);

	delay6 : component alt_dspbuilder_delay_GNALDIUCHM
		generic map (
			ClockPhase => "1",
			BitPattern => "000000000001",
			width      => 12,
			use_init   => 0,
			delay      => 6
		)
		port map (
			input  => logical_bus_operator3_result_wire, --      input.wire
			clock  => clock_0_clock_output_clk,          -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,        --           .reset
			output => delay6_output_wire,                --     output.wire
			sclr   => delay6sclrgnd_output_wire,         --       sclr.wire
			ena    => clken_0_output_wire                --        ena.wire
		);

	delay6sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delay6sclrgnd_output_wire  -- output.wire
		);

	delay5 : component alt_dspbuilder_delay_GNSPCBEWTM
		generic map (
			ClockPhase => "1",
			BitPattern => "0000000001",
			width      => 10,
			use_init   => 0,
			delay      => 6
		)
		port map (
			input  => logical_bus_operator2_result_wire, --      input.wire
			clock  => clock_0_clock_output_clk,          -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,        --           .reset
			output => delay5_output_wire,                --     output.wire
			sclr   => delay5sclrgnd_output_wire,         --       sclr.wire
			ena    => clken_0_output_wire                --        ena.wire
		);

	delay5sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delay5sclrgnd_output_wire  -- output.wire
		);

	memory_delay : component alt_dspbuilder_memdelay_GNOQUXON7R
		generic map (
			RAMTYPE => "AUTO",
			WIDTH   => 8,
			DELAY   => 27
		)
		port map (
			clock     => clock_0_clock_output_clk,             -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,           --           .reset
			input     => data_22_0_output_wire,                --      input.wire
			output    => memory_delay_output_wire,             --     output.wire
			user_aclr => memory_delayuser_aclrgnd_output_wire, --  user_aclr.wire
			ena       => clken_0_output_wire                   --        ena.wire
		);

	memory_delayuser_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => memory_delayuser_aclrgnd_output_wire  -- output.wire
		);

	delay4 : component alt_dspbuilder_delay_GNMDMEZDYK
		generic map (
			ClockPhase => "1",
			BitPattern => "00000001",
			width      => 8,
			use_init   => 0,
			delay      => 6
		)
		port map (
			input  => data_04_0_output_wire,      --      input.wire
			clock  => clock_0_clock_output_clk,   -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset, --           .reset
			output => delay4_output_wire,         --     output.wire
			sclr   => delay4sclrgnd_output_wire,  --       sclr.wire
			ena    => clken_0_output_wire         --        ena.wire
		);

	delay4sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delay4sclrgnd_output_wire  -- output.wire
		);

	delay3 : component alt_dspbuilder_delay_GNSPCBEWTM
		generic map (
			ClockPhase => "1",
			BitPattern => "0000000001",
			width      => 10,
			use_init   => 0,
			delay      => 6
		)
		port map (
			input  => logical_bus_operator1_result_wire, --      input.wire
			clock  => clock_0_clock_output_clk,          -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,        --           .reset
			output => delay3_output_wire,                --     output.wire
			sclr   => delay3sclrgnd_output_wire,         --       sclr.wire
			ena    => clken_0_output_wire                --        ena.wire
		);

	delay3sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delay3sclrgnd_output_wire  -- output.wire
		);

	delay9 : component alt_dspbuilder_delay_GNSPCBEWTM
		generic map (
			ClockPhase => "1",
			BitPattern => "0000000001",
			width      => 10,
			use_init   => 0,
			delay      => 6
		)
		port map (
			input  => logical_bus_operator5_result_wire, --      input.wire
			clock  => clock_0_clock_output_clk,          -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,        --           .reset
			output => delay9_output_wire,                --     output.wire
			sclr   => delay9sclrgnd_output_wire,         --       sclr.wire
			ena    => clken_0_output_wire                --        ena.wire
		);

	delay9sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delay9sclrgnd_output_wire  -- output.wire
		);

	delay8 : component alt_dspbuilder_delay_GNALDIUCHM
		generic map (
			ClockPhase => "1",
			BitPattern => "000000000001",
			width      => 12,
			use_init   => 0,
			delay      => 6
		)
		port map (
			input  => logical_bus_operator4_result_wire, --      input.wire
			clock  => clock_0_clock_output_clk,          -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,        --           .reset
			output => delay8_output_wire,                --     output.wire
			sclr   => delay8sclrgnd_output_wire,         --       sclr.wire
			ena    => clken_0_output_wire                --        ena.wire
		);

	delay8sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delay8sclrgnd_output_wire  -- output.wire
		);

	delay7 : component alt_dspbuilder_delay_GN2KYXQF4S
		generic map (
			ClockPhase => "1",
			BitPattern => "000000000000001",
			width      => 15,
			use_init   => 0,
			delay      => 1
		)
		port map (
			input  => gain1_output_wire,          --      input.wire
			clock  => clock_0_clock_output_clk,   -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset, --           .reset
			output => delay7_output_wire,         --     output.wire
			sclr   => delay7sclrgnd_output_wire,  --       sclr.wire
			ena    => clken_0_output_wire         --        ena.wire
		);

	delay7sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delay7sclrgnd_output_wire  -- output.wire
		);

	cast133 : component alt_dspbuilder_cast_GNUW2C7J4Q
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => data_02_0_output_wire, --  input.wire
			output => cast133_output_wire    -- output.wire
		);

	cast134 : component alt_dspbuilder_cast_GNUW2C7J4Q
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => data_12_0_output_wire, --  input.wire
			output => cast134_output_wire    -- output.wire
		);

	cast135 : component alt_dspbuilder_cast_GNUW2C7J4Q
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => data_20_0_output_wire, --  input.wire
			output => cast135_output_wire    -- output.wire
		);

	cast136 : component alt_dspbuilder_cast_GNUW2C7J4Q
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => data_21_0_output_wire, --  input.wire
			output => cast136_output_wire    -- output.wire
		);

	cast137 : component alt_dspbuilder_cast_GNUW2C7J4Q
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => data_22_0_output_wire, --  input.wire
			output => cast137_output_wire    -- output.wire
		);

	cast138 : component alt_dspbuilder_cast_GNUW2C7J4Q
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => data_23_0_output_wire, --  input.wire
			output => cast138_output_wire    -- output.wire
		);

	cast139 : component alt_dspbuilder_cast_GNUW2C7J4Q
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => data_24_0_output_wire, --  input.wire
			output => cast139_output_wire    -- output.wire
		);

	cast140 : component alt_dspbuilder_cast_GNUW2C7J4Q
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => data_32_0_output_wire, --  input.wire
			output => cast140_output_wire    -- output.wire
		);

	cast141 : component alt_dspbuilder_cast_GNUW2C7J4Q
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => data_42_0_output_wire, --  input.wire
			output => cast141_output_wire    -- output.wire
		);

	cast142 : component alt_dspbuilder_cast_GNNDZ2WJEB
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => data_01_0_output_wire, --  input.wire
			output => cast142_output_wire    -- output.wire
		);

	cast143 : component alt_dspbuilder_cast_GNNDZ2WJEB
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => data_03_0_output_wire, --  input.wire
			output => cast143_output_wire    -- output.wire
		);

	cast144 : component alt_dspbuilder_cast_GNNDZ2WJEB
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => data_41_0_output_wire, --  input.wire
			output => cast144_output_wire    -- output.wire
		);

	cast145 : component alt_dspbuilder_cast_GNNDZ2WJEB
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => data_43_0_output_wire, --  input.wire
			output => cast145_output_wire    -- output.wire
		);

	cast146 : component alt_dspbuilder_cast_GNNDZ2WJEB
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => data_10_0_output_wire, --  input.wire
			output => cast146_output_wire    -- output.wire
		);

	cast147 : component alt_dspbuilder_cast_GNUJN4ENCM
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => data_11_0_output_wire, --  input.wire
			output => cast147_output_wire    -- output.wire
		);

	cast148 : component alt_dspbuilder_cast_GNUJN4ENCM
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => data_13_0_output_wire, --  input.wire
			output => cast148_output_wire    -- output.wire
		);

	cast149 : component alt_dspbuilder_cast_GNNDZ2WJEB
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => data_14_0_output_wire, --  input.wire
			output => cast149_output_wire    -- output.wire
		);

	cast150 : component alt_dspbuilder_cast_GNNDZ2WJEB
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => data_30_0_output_wire, --  input.wire
			output => cast150_output_wire    -- output.wire
		);

	cast151 : component alt_dspbuilder_cast_GNUJN4ENCM
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => data_31_0_output_wire, --  input.wire
			output => cast151_output_wire    -- output.wire
		);

	cast152 : component alt_dspbuilder_cast_GNUJN4ENCM
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => data_33_0_output_wire, --  input.wire
			output => cast152_output_wire    -- output.wire
		);

	cast153 : component alt_dspbuilder_cast_GNNDZ2WJEB
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => data_34_0_output_wire, --  input.wire
			output => cast153_output_wire    -- output.wire
		);

	cast154 : component alt_dspbuilder_cast_GNBZR5PMEK
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => memory_delay_output_wire, --  input.wire
			output => cast154_output_wire       -- output.wire
		);

	cast155 : component alt_dspbuilder_cast_GN4Q52ZVBU
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => parallel_adder_subtractor_result_wire, --  input.wire
			output => cast155_output_wire                    -- output.wire
		);

	cast156 : component alt_dspbuilder_cast_GNT75CKW5G
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => delay_output_wire,   --  input.wire
			output => cast156_output_wire  -- output.wire
		);

	cast157 : component alt_dspbuilder_cast_GNSGOYMYTM
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => delay1_output_wire,  --  input.wire
			output => cast157_output_wire  -- output.wire
		);

	cast158 : component alt_dspbuilder_cast_GNYETX3347
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => delay2_output_wire,  --  input.wire
			output => cast158_output_wire  -- output.wire
		);

	cast159 : component alt_dspbuilder_cast_GNSGOYMYTM
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => delay3_output_wire,  --  input.wire
			output => cast159_output_wire  -- output.wire
		);

	cast160 : component alt_dspbuilder_cast_GNT75CKW5G
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => delay4_output_wire,  --  input.wire
			output => cast160_output_wire  -- output.wire
		);

	cast161 : component alt_dspbuilder_cast_GNSGOYMYTM
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => delay5_output_wire,  --  input.wire
			output => cast161_output_wire  -- output.wire
		);

	cast162 : component alt_dspbuilder_cast_GNPGJSMS3Z
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => delay6_output_wire,  --  input.wire
			output => cast162_output_wire  -- output.wire
		);

	cast163 : component alt_dspbuilder_cast_GNZCDPTGZG
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => delay7_output_wire,  --  input.wire
			output => cast163_output_wire  -- output.wire
		);

	cast164 : component alt_dspbuilder_cast_GNPGJSMS3Z
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => delay8_output_wire,  --  input.wire
			output => cast164_output_wire  -- output.wire
		);

	cast165 : component alt_dspbuilder_cast_GNSGOYMYTM
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => delay9_output_wire,  --  input.wire
			output => cast165_output_wire  -- output.wire
		);

	cast166 : component alt_dspbuilder_cast_GNYETX3347
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => delay10_output_wire, --  input.wire
			output => cast166_output_wire  -- output.wire
		);

	cast167 : component alt_dspbuilder_cast_GNZCDPTGZG
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => delay11_output_wire, --  input.wire
			output => cast167_output_wire  -- output.wire
		);

	cast168 : component alt_dspbuilder_cast_GNZCDPTGZG
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => delay13_output_wire, --  input.wire
			output => cast168_output_wire  -- output.wire
		);

	cast169 : component alt_dspbuilder_cast_GNYETX3347
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => delay14_output_wire, --  input.wire
			output => cast169_output_wire  -- output.wire
		);

	cast170 : component alt_dspbuilder_cast_GNSGOYMYTM
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => delay12_output_wire, --  input.wire
			output => cast170_output_wire  -- output.wire
		);

	cast171 : component alt_dspbuilder_cast_GNPGJSMS3Z
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => delay15_output_wire, --  input.wire
			output => cast171_output_wire  -- output.wire
		);

	cast172 : component alt_dspbuilder_cast_GNZCDPTGZG
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => delay16_output_wire, --  input.wire
			output => cast172_output_wire  -- output.wire
		);

	cast173 : component alt_dspbuilder_cast_GNPGJSMS3Z
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => delay17_output_wire, --  input.wire
			output => cast173_output_wire  -- output.wire
		);

	cast174 : component alt_dspbuilder_cast_GNSGOYMYTM
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => delay18_output_wire, --  input.wire
			output => cast174_output_wire  -- output.wire
		);

	cast175 : component alt_dspbuilder_cast_GNT75CKW5G
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => delay19_output_wire, --  input.wire
			output => cast175_output_wire  -- output.wire
		);

	cast176 : component alt_dspbuilder_cast_GNSGOYMYTM
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => delay20_output_wire, --  input.wire
			output => cast176_output_wire  -- output.wire
		);

	cast177 : component alt_dspbuilder_cast_GNYETX3347
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => delay21_output_wire, --  input.wire
			output => cast177_output_wire  -- output.wire
		);

	cast178 : component alt_dspbuilder_cast_GNSGOYMYTM
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => delay22_output_wire, --  input.wire
			output => cast178_output_wire  -- output.wire
		);

	cast179 : component alt_dspbuilder_cast_GNT75CKW5G
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => delay23_output_wire, --  input.wire
			output => cast179_output_wire  -- output.wire
		);

	cast180 : component alt_dspbuilder_cast_GNBZR5PMEK
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => round_dataout_wire,  --  input.wire
			output => cast180_output_wire  -- output.wire
		);

end architecture rtl; -- of gaussian_ip_GN_gaussian_ip_Fusion_Decomposition_2_multiplier_accumulator
