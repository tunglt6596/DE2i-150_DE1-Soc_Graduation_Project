-- localedgepreserve_GN_localedgepreserve_Fusion.vhd

-- Generated using ACDS version 17.1 590

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity localedgepreserve_GN_localedgepreserve_Fusion is
	port (
		eof_in    : in  std_logic                    := '0';             --    eof_in.wire
		valid_out : out std_logic;                                       -- valid_out.wire
		pixel_in  : in  std_logic_vector(7 downto 0) := (others => '0'); --  pixel_in.wire
		valid1_in : in  std_logic                    := '0';             -- valid1_in.wire
		eof2_in   : in  std_logic                    := '0';             --   eof2_in.wire
		Clock     : in  std_logic                    := '0';             --     Clock.clk
		reset     : in  std_logic                    := '0';             --          .reset
		pixel1_in : in  std_logic_vector(7 downto 0) := (others => '0'); -- pixel1_in.wire
		sof_out   : out std_logic;                                       --   sof_out.wire
		eof1_in   : in  std_logic                    := '0';             --   eof1_in.wire
		eof_out   : out std_logic;                                       --   eof_out.wire
		pixel2_in : in  std_logic_vector(7 downto 0) := (others => '0'); -- pixel2_in.wire
		pixel_out : out std_logic_vector(8 downto 0);                    -- pixel_out.wire
		valid2_in : in  std_logic                    := '0';             -- valid2_in.wire
		valid_in  : in  std_logic                    := '0'              --  valid_in.wire
	);
end entity localedgepreserve_GN_localedgepreserve_Fusion;

architecture rtl of localedgepreserve_GN_localedgepreserve_Fusion is
	component alt_dspbuilder_clock_GNQFU4PUDH is
		port (
			aclr      : in  std_logic := 'X'; -- reset
			aclr_n    : in  std_logic := 'X'; -- reset_n
			aclr_out  : out std_logic;        -- reset
			clock     : in  std_logic := 'X'; -- clk
			clock_out : out std_logic         -- clk
		);
	end component alt_dspbuilder_clock_GNQFU4PUDH;

	component alt_dspbuilder_port_GN37ALZBS4 is
		port (
			input  : in  std_logic := 'X'; -- wire
			output : out std_logic         -- wire
		);
	end component alt_dspbuilder_port_GN37ALZBS4;

	component alt_dspbuilder_multiplier_GNSFKO7633 is
		generic (
			aWidth                         : natural := 8;
			Signed                         : natural := 0;
			bWidth                         : natural := 8;
			DEDICATED_MULTIPLIER_CIRCUITRY : string  := "AUTO";
			pipeline                       : integer := 0;
			OutputLsb                      : integer := 0;
			OutputMsb                      : integer := 8
		);
		port (
			aclr      : in  std_logic                                          := 'X';             -- clk
			clock     : in  std_logic                                          := 'X';             -- clk
			dataa     : in  std_logic_vector(aWidth-1 downto 0)                := (others => 'X'); -- wire
			datab     : in  std_logic_vector(bWidth-1 downto 0)                := (others => 'X'); -- wire
			ena       : in  std_logic                                          := 'X';             -- wire
			result    : out std_logic_vector(OutputMsb-OutputLsb+1-1 downto 0);                    -- wire
			user_aclr : in  std_logic                                          := 'X'              -- wire
		);
	end component alt_dspbuilder_multiplier_GNSFKO7633;

	component alt_dspbuilder_gnd_GN is
		port (
			output : out std_logic   -- wire
		);
	end component alt_dspbuilder_gnd_GN;

	component alt_dspbuilder_cast_GNUYRTQ4QH is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(23 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNUYRTQ4QH;

	component alt_dspbuilder_multiplexer_GNIM5IEXF4 is
		generic (
			number_inputs          : natural  := 4;
			pipeline               : natural  := 0;
			width                  : positive := 8;
			HDLTYPE                : string   := "STD_LOGIC_VECTOR";
			use_one_hot_select_bus : natural  := 0
		);
		port (
			clock     : in  std_logic                    := 'X';             -- clk
			aclr      : in  std_logic                    := 'X';             -- reset
			sel       : in  std_logic_vector(0 downto 0) := (others => 'X'); -- wire
			result    : out std_logic_vector(8 downto 0);                    -- wire
			ena       : in  std_logic                    := 'X';             -- wire
			user_aclr : in  std_logic                    := 'X';             -- wire
			in0       : in  std_logic_vector(8 downto 0) := (others => 'X'); -- wire
			in1       : in  std_logic_vector(8 downto 0) := (others => 'X')  -- wire
		);
	end component alt_dspbuilder_multiplexer_GNIM5IEXF4;

	component alt_dspbuilder_vcc_GN is
		port (
			output : out std_logic   -- wire
		);
	end component alt_dspbuilder_vcc_GN;

	component alt_dspbuilder_port_GNA5S4SQDN is
		port (
			input  : in  std_logic_vector(7 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(7 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNA5S4SQDN;

	component localedgepreserve_GN_localedgepreserve_Fusion_Cal_Image_Out_2 is
		port (
			pixel_in : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- wire
			a_in     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- wire
			b_in     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- wire
			ir       : out std_logic_vector(7 downto 0);                     -- wire
			p_ir     : out std_logic_vector(15 downto 0);                    -- wire
			Clock    : in  std_logic                     := 'X';             -- clk
			reset    : in  std_logic                     := 'X';             -- reset
			valid_in : in  std_logic                     := 'X'              -- wire
		);
	end component localedgepreserve_GN_localedgepreserve_Fusion_Cal_Image_Out_2;

	component alt_dspbuilder_delay_GNCY3KEQXH is
		generic (
			ClockPhase : string   := "1";
			BitPattern : string   := "00000001";
			width      : positive := 8;
			use_init   : natural  := 0;
			delay      : positive := 1
		);
		port (
			aclr   : in  std_logic                          := 'X';             -- clk
			clock  : in  std_logic                          := 'X';             -- clk
			ena    : in  std_logic                          := 'X';             -- wire
			input  : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(width-1 downto 0);                    -- wire
			sclr   : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_delay_GNCY3KEQXH;

	component localedgepreserve_GN_localedgepreserve_Fusion_Cal_Image_Out_1 is
		port (
			valid_in : in  std_logic                     := 'X';             -- wire
			p_vis    : out std_logic_vector(15 downto 0);                    -- wire
			a_in     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- wire
			pixel_in : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- wire
			Clock    : in  std_logic                     := 'X';             -- clk
			reset    : in  std_logic                     := 'X';             -- reset
			b_in     : in  std_logic_vector(15 downto 0) := (others => 'X')  -- wire
		);
	end component localedgepreserve_GN_localedgepreserve_Fusion_Cal_Image_Out_1;

	component alt_dspbuilder_comparator_GN is
		generic (
			Operator  : string  := "Altaeb";
			lpm_width : natural := 8
		);
		port (
			clock  : in  std_logic                              := 'X';             -- clk
			dataa  : in  std_logic_vector(lpm_width-1 downto 0) := (others => 'X'); -- wire
			datab  : in  std_logic_vector(lpm_width-1 downto 0) := (others => 'X'); -- wire
			result : out std_logic;                                                 -- wire
			sclr   : in  std_logic                              := 'X'              -- clk
		);
	end component alt_dspbuilder_comparator_GN;

	component localedgepreserve_GN_localedgepreserve_Fusion_generate_signals is
		port (
			eof_in    : in  std_logic := 'X'; -- wire
			sof_out   : out std_logic;        -- wire
			valid_in  : in  std_logic := 'X'; -- wire
			valid_out : out std_logic;        -- wire
			Clock     : in  std_logic := 'X'; -- clk
			reset     : in  std_logic := 'X'; -- reset
			eof_out   : out std_logic         -- wire
		);
	end component localedgepreserve_GN_localedgepreserve_Fusion_generate_signals;

	component alt_dspbuilder_pipelined_adder_GNTWZRTG4I is
		generic (
			pipeline : integer := 0;
			width    : natural := 0
		);
		port (
			aclr      : in  std_logic                          := 'X';             -- clk
			add_sub   : in  std_logic                          := 'X';             -- wire
			cin       : in  std_logic                          := 'X';             -- wire
			clock     : in  std_logic                          := 'X';             -- clk
			cout      : out std_logic;                                             -- wire
			dataa     : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			datab     : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			ena       : in  std_logic                          := 'X';             -- wire
			result    : out std_logic_vector(width-1 downto 0);                    -- wire
			user_aclr : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_pipelined_adder_GNTWZRTG4I;

	component alt_dspbuilder_cast_GNEBWH7Z3U is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(23 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNEBWH7Z3U;

	component alt_dspbuilder_cast_GN7IYG3D6O is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(24 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(8 downto 0)                      -- wire
		);
	end component alt_dspbuilder_cast_GN7IYG3D6O;

	component alt_dspbuilder_cast_GNEL6FJM3V is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(16 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNEL6FJM3V;

	component alt_dspbuilder_constant_GNSVSRQZMI is
		generic (
			BitPattern : string  := "0000";
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(7 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GNSVSRQZMI;

	component alt_dspbuilder_constant_GNQQLU6SNF is
		generic (
			BitPattern : string  := "0000";
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(16 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GNQQLU6SNF;

	component alt_dspbuilder_constant_GNP7U2HOAO is
		generic (
			BitPattern : string  := "0000";
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(8 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GNP7U2HOAO;

	component alt_dspbuilder_bus_concat_GNU3KBQ5HN is
		generic (
			widthA : natural := 8;
			widthB : natural := 8
		);
		port (
			a      : in  std_logic_vector(widthA-1 downto 0)        := (others => 'X'); -- wire
			aclr   : in  std_logic                                  := 'X';             -- clk
			b      : in  std_logic_vector(widthB-1 downto 0)        := (others => 'X'); -- wire
			clock  : in  std_logic                                  := 'X';             -- clk
			output : out std_logic_vector(widthA+widthB-1 downto 0)                     -- wire
		);
	end component alt_dspbuilder_bus_concat_GNU3KBQ5HN;

	component alt_dspbuilder_bus_concat_GN7K3OAUCY is
		generic (
			widthA : natural := 8;
			widthB : natural := 8
		);
		port (
			a      : in  std_logic_vector(widthA-1 downto 0)        := (others => 'X'); -- wire
			aclr   : in  std_logic                                  := 'X';             -- clk
			b      : in  std_logic_vector(widthB-1 downto 0)        := (others => 'X'); -- wire
			clock  : in  std_logic                                  := 'X';             -- clk
			output : out std_logic_vector(widthA+widthB-1 downto 0)                     -- wire
		);
	end component alt_dspbuilder_bus_concat_GN7K3OAUCY;

	component alt_dspbuilder_constant_GNCWI5QDAD is
		generic (
			BitPattern : string  := "0000";
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(15 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GNCWI5QDAD;

	component alt_dspbuilder_constant_GNC5NOVIJT is
		generic (
			BitPattern : string  := "0000";
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(7 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GNC5NOVIJT;

	component alt_dspbuilder_constant_GNDEA2MM7Q is
		generic (
			BitPattern : string  := "0000";
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(16 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GNDEA2MM7Q;

	component alt_dspbuilder_port_GNJVFJM3AT is
		port (
			input  : in  std_logic_vector(8 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(8 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNJVFJM3AT;

	component alt_dspbuilder_multiplexer_GNMRY6PWYH is
		generic (
			number_inputs          : natural  := 4;
			pipeline               : natural  := 0;
			width                  : positive := 8;
			HDLTYPE                : string   := "STD_LOGIC_VECTOR";
			use_one_hot_select_bus : natural  := 0
		);
		port (
			clock     : in  std_logic                     := 'X';             -- clk
			aclr      : in  std_logic                     := 'X';             -- reset
			sel       : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- wire
			result    : out std_logic_vector(16 downto 0);                    -- wire
			ena       : in  std_logic                     := 'X';             -- wire
			user_aclr : in  std_logic                     := 'X';             -- wire
			in0       : in  std_logic_vector(16 downto 0) := (others => 'X'); -- wire
			in1       : in  std_logic_vector(16 downto 0) := (others => 'X')  -- wire
		);
	end component alt_dspbuilder_multiplexer_GNMRY6PWYH;

	component localedgepreserve_GN_localedgepreserve_Fusion_Cal_A_B_2 is
		port (
			eof_in    : in  std_logic                     := 'X';             -- wire
			a_out     : out std_logic_vector(15 downto 0);                    -- wire
			pixel_in  : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- wire
			b_out     : out std_logic_vector(15 downto 0);                    -- wire
			pixel_out : out std_logic_vector(7 downto 0);                     -- wire
			Clock     : in  std_logic                     := 'X';             -- clk
			reset     : in  std_logic                     := 'X';             -- reset
			grad_in   : in  std_logic_vector(10 downto 0) := (others => 'X'); -- wire
			eof_out   : out std_logic;                                        -- wire
			valid_in  : in  std_logic                     := 'X';             -- wire
			valid_out : out std_logic                                         -- wire
		);
	end component localedgepreserve_GN_localedgepreserve_Fusion_Cal_A_B_2;

	component alt_dspbuilder_pipelined_adder_GNWEIMU3MK is
		generic (
			pipeline : integer := 0;
			width    : natural := 0
		);
		port (
			aclr      : in  std_logic                          := 'X';             -- clk
			add_sub   : in  std_logic                          := 'X';             -- wire
			cin       : in  std_logic                          := 'X';             -- wire
			clock     : in  std_logic                          := 'X';             -- clk
			cout      : out std_logic;                                             -- wire
			dataa     : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			datab     : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			ena       : in  std_logic                          := 'X';             -- wire
			result    : out std_logic_vector(width-1 downto 0);                    -- wire
			user_aclr : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_pipelined_adder_GNWEIMU3MK;

	component localedgepreserve_GN_localedgepreserve_Fusion_Cal_A_B_1 is
		port (
			eof_in    : in  std_logic                     := 'X';             -- wire
			b_out     : out std_logic_vector(15 downto 0);                    -- wire
			valid_out : out std_logic;                                        -- wire
			a_out     : out std_logic_vector(15 downto 0);                    -- wire
			pixel_out : out std_logic_vector(7 downto 0);                     -- wire
			grad_in   : in  std_logic_vector(10 downto 0) := (others => 'X'); -- wire
			valid_in  : in  std_logic                     := 'X';             -- wire
			pixel_in  : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- wire
			Clock     : in  std_logic                     := 'X';             -- clk
			reset     : in  std_logic                     := 'X'              -- reset
		);
	end component localedgepreserve_GN_localedgepreserve_Fusion_Cal_A_B_1;

	component alt_dspbuilder_memdelay_GNBRIKDQTV is
		generic (
			RAMTYPE : string   := "AUTO";
			WIDTH   : positive := 8;
			DELAY   : positive := 1
		);
		port (
			aclr      : in  std_logic                          := 'X';             -- clk
			clock     : in  std_logic                          := 'X';             -- clk
			ena       : in  std_logic                          := 'X';             -- wire
			input     : in  std_logic_vector(WIDTH-1 downto 0) := (others => 'X'); -- wire
			output    : out std_logic_vector(WIDTH-1 downto 0);                    -- wire
			user_aclr : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_memdelay_GNBRIKDQTV;

	component alt_dspbuilder_delay_GNIDQK4WDH is
		generic (
			ClockPhase : string   := "1";
			BitPattern : string   := "00000001";
			width      : positive := 8;
			use_init   : natural  := 0;
			delay      : positive := 1
		);
		port (
			aclr   : in  std_logic                          := 'X';             -- clk
			clock  : in  std_logic                          := 'X';             -- clk
			ena    : in  std_logic                          := 'X';             -- wire
			input  : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(width-1 downto 0);                    -- wire
			sclr   : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_delay_GNIDQK4WDH;

	component localedgepreserve_GN_localedgepreserve_Fusion_Cal_Weight is
		port (
			max_out   : out std_logic_vector(31 downto 0);                    -- wire
			pixel_in  : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- wire
			eof_in    : in  std_logic                     := 'X';             -- wire
			valid_in  : in  std_logic                     := 'X';             -- wire
			value_out : out std_logic_vector(31 downto 0);                    -- wire
			Clock     : in  std_logic                     := 'X';             -- clk
			reset     : in  std_logic                     := 'X';             -- reset
			addr_in   : in  std_logic_vector(7 downto 0)  := (others => 'X')  -- wire
		);
	end component localedgepreserve_GN_localedgepreserve_Fusion_Cal_Weight;

	component localedgepreserve_GN_localedgepreserve_Fusion_Cal_Magnitude_Gradient_2 is
		port (
			sof_out   : out std_logic;                                        -- wire
			pixel_out : out std_logic_vector(7 downto 0);                     -- wire
			eof_out   : out std_logic;                                        -- wire
			pixel_in  : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- wire
			grad_out  : out std_logic_vector(10 downto 0);                    -- wire
			valid_out : out std_logic;                                        -- wire
			valid_in  : in  std_logic                     := 'X';             -- wire
			Clock     : in  std_logic                     := 'X';             -- clk
			reset     : in  std_logic                     := 'X';             -- reset
			eof_in    : in  std_logic                     := 'X'              -- wire
		);
	end component localedgepreserve_GN_localedgepreserve_Fusion_Cal_Magnitude_Gradient_2;

	component localedgepreserve_GN_localedgepreserve_Fusion_Cal_Magnitude_Gradient_1 is
		port (
			eof_in    : in  std_logic                     := 'X';             -- wire
			grad_out  : out std_logic_vector(10 downto 0);                    -- wire
			pixel_out : out std_logic_vector(7 downto 0);                     -- wire
			valid_in  : in  std_logic                     := 'X';             -- wire
			eof_out   : out std_logic;                                        -- wire
			Clock     : in  std_logic                     := 'X';             -- clk
			reset     : in  std_logic                     := 'X';             -- reset
			pixel_in  : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- wire
			valid_out : out std_logic                                         -- wire
		);
	end component localedgepreserve_GN_localedgepreserve_Fusion_Cal_Magnitude_Gradient_1;

	component alt_dspbuilder_memdelay_GN3YPLAG7W is
		generic (
			RAMTYPE : string   := "AUTO";
			WIDTH   : positive := 8;
			DELAY   : positive := 1
		);
		port (
			aclr      : in  std_logic                          := 'X';             -- clk
			clock     : in  std_logic                          := 'X';             -- clk
			ena       : in  std_logic                          := 'X';             -- wire
			input     : in  std_logic_vector(WIDTH-1 downto 0) := (others => 'X'); -- wire
			output    : out std_logic_vector(WIDTH-1 downto 0);                    -- wire
			user_aclr : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_memdelay_GN3YPLAG7W;

	component div is
		port (
			clk : in  std_logic                     := 'X';             -- clk
			d   : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			ena : in  std_logic                     := 'X';             -- wire
			q   : out std_logic_vector(23 downto 0);                    -- wire
			z   : in  std_logic_vector(47 downto 0) := (others => 'X')  -- wire
		);
	end component div;

	component alt_dspbuilder_cast_GNA5TAMWCZ is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(23 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNA5TAMWCZ;

	component alt_dspbuilder_cast_GNPFJ7B3O7 is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(8 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(9 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNPFJ7B3O7;

	component alt_dspbuilder_cast_GN7YNIFSF6 is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(16 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(17 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GN7YNIFSF6;

	component alt_dspbuilder_cast_GNKD3JEUSD is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(47 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(47 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNKD3JEUSD;

	component alt_dspbuilder_cast_GN5P6ORZXA is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(23 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GN5P6ORZXA;

	component alt_dspbuilder_cast_GNEIIG67TZ is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(23 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNEIIG67TZ;

	component alt_dspbuilder_cast_GN46N4UJ5S is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic                    := 'X'; -- wire
			output : out std_logic_vector(0 downto 0)         -- wire
		);
	end component alt_dspbuilder_cast_GN46N4UJ5S;

	component alt_dspbuilder_cast_GNXDXNUGW4 is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(7 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(8 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNXDXNUGW4;

	component alt_dspbuilder_cast_GNJ6DWMNK6 is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(24 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNJ6DWMNK6;

	signal multiplier1user_aclrgnd_output_wire                                : std_logic;                     -- Multiplier1user_aclrGND:output -> Multiplier1:user_aclr
	signal multiplexeruser_aclrgnd_output_wire                                : std_logic;                     -- Multiplexeruser_aclrGND:output -> Multiplexer:user_aclr
	signal multiplexerenavcc_output_wire                                      : std_logic;                     -- MultiplexerenaVCC:output -> Multiplexer:ena
	signal delaysclrgnd_output_wire                                           : std_logic;                     -- DelaysclrGND:output -> Delay:sclr
	signal pipelined_adder1user_aclrgnd_output_wire                           : std_logic;                     -- Pipelined_Adder1user_aclrGND:output -> Pipelined_Adder1:user_aclr
	signal multiplexer1user_aclrgnd_output_wire                               : std_logic;                     -- Multiplexer1user_aclrGND:output -> Multiplexer1:user_aclr
	signal multiplexer1enavcc_output_wire                                     : std_logic;                     -- Multiplexer1enaVCC:output -> Multiplexer1:ena
	signal pipelined_adderuser_aclrgnd_output_wire                            : std_logic;                     -- Pipelined_Adderuser_aclrGND:output -> Pipelined_Adder:user_aclr
	signal memory_delay1user_aclrgnd_output_wire                              : std_logic;                     -- Memory_Delay1user_aclrGND:output -> Memory_Delay1:user_aclr
	signal multiplieruser_aclrgnd_output_wire                                 : std_logic;                     -- Multiplieruser_aclrGND:output -> Multiplier:user_aclr
	signal delay1sclrgnd_output_wire                                          : std_logic;                     -- Delay1sclrGND:output -> Delay1:sclr
	signal memory_delayuser_aclrgnd_output_wire                               : std_logic;                     -- Memory_Delayuser_aclrGND:output -> Memory_Delay:user_aclr
	signal bus_concatenation2_output_wire                                     : std_logic_vector(39 downto 0); -- Bus_Concatenation2:output -> Bus_Concatenation3:b
	signal binary_point_casting1_output_wire                                  : std_logic_vector(23 downto 0); -- Binary_Point_Casting1:output -> Bus_Conversion1:input
	signal bus_conversion2_output_wire                                        : std_logic_vector(23 downto 0); -- Bus_Conversion2:output -> Binary_Point_Casting3:input
	signal bus_conversion3_output_wire                                        : std_logic_vector(23 downto 0); -- Bus_Conversion3:output -> Binary_Point_Casting2:input
	signal constant6_output_wire                                              : std_logic_vector(15 downto 0); -- Constant6:output -> Bus_Concatenation2:b
	signal constant7_output_wire                                              : std_logic_vector(7 downto 0);  -- Constant7:output -> Bus_Concatenation3:a
	signal bus_conversion1_output_wire                                        : std_logic_vector(16 downto 0); -- Bus_Conversion1:output -> [Delay1:input, Multiplier:dataa, Pipelined_Adder:datab]
	signal localedgepreserve_fusion_cal_magnitude_gradient_2_0_pixel_out_wire : std_logic_vector(7 downto 0);  -- localedgepreserve_Fusion_Cal_Magnitude_Gradient_2_0:pixel_out -> localedgepreserve_Fusion_Cal_A_B_2_0:pixel_in
	signal localedgepreserve_fusion_cal_magnitude_gradient_2_0_grad_out_wire  : std_logic_vector(10 downto 0); -- localedgepreserve_Fusion_Cal_Magnitude_Gradient_2_0:grad_out -> localedgepreserve_Fusion_Cal_A_B_2_0:grad_in
	signal localedgepreserve_fusion_cal_a_b_2_0_pixel_out_wire                : std_logic_vector(7 downto 0);  -- localedgepreserve_Fusion_Cal_A_B_2_0:pixel_out -> localedgepreserve_Fusion_Cal_Image_Out_2_0:pixel_in
	signal pixel2_in_0_output_wire                                            : std_logic_vector(7 downto 0);  -- pixel2_in_0:output -> localedgepreserve_Fusion_Cal_Magnitude_Gradient_2_0:pixel_in
	signal valid2_in_0_output_wire                                            : std_logic;                     -- valid2_in_0:output -> localedgepreserve_Fusion_Cal_Magnitude_Gradient_2_0:valid_in
	signal eof2_in_0_output_wire                                              : std_logic;                     -- eof2_in_0:output -> localedgepreserve_Fusion_Cal_Magnitude_Gradient_2_0:eof_in
	signal localedgepreserve_fusion_cal_magnitude_gradient_1_0_pixel_out_wire : std_logic_vector(7 downto 0);  -- localedgepreserve_Fusion_Cal_Magnitude_Gradient_1_0:pixel_out -> localedgepreserve_Fusion_Cal_A_B_1_0:pixel_in
	signal localedgepreserve_fusion_cal_a_b_2_0_a_out_wire                    : std_logic_vector(15 downto 0); -- localedgepreserve_Fusion_Cal_A_B_2_0:a_out -> localedgepreserve_Fusion_Cal_Image_Out_2_0:a_in
	signal localedgepreserve_fusion_cal_magnitude_gradient_1_0_grad_out_wire  : std_logic_vector(10 downto 0); -- localedgepreserve_Fusion_Cal_Magnitude_Gradient_1_0:grad_out -> localedgepreserve_Fusion_Cal_A_B_1_0:grad_in
	signal localedgepreserve_fusion_cal_a_b_1_0_pixel_out_wire                : std_logic_vector(7 downto 0);  -- localedgepreserve_Fusion_Cal_A_B_1_0:pixel_out -> localedgepreserve_Fusion_Cal_Image_Out_1_0:pixel_in
	signal pixel1_in_0_output_wire                                            : std_logic_vector(7 downto 0);  -- pixel1_in_0:output -> localedgepreserve_Fusion_Cal_Magnitude_Gradient_1_0:pixel_in
	signal localedgepreserve_fusion_cal_a_b_2_0_valid_out_wire                : std_logic;                     -- localedgepreserve_Fusion_Cal_A_B_2_0:valid_out -> [Delay1:ena, Delay:ena, Divider:ena, Memory_Delay1:ena, Memory_Delay:ena, Multiplier1:ena, Multiplier:ena, Pipelined_Adder1:ena, Pipelined_Adder:ena, localedgepreserve_Fusion_Cal_Image_Out_2_0:valid_in, localedgepreserve_Fusion_generate_signals_0:valid_in]
	signal localedgepreserve_fusion_cal_weight_0_max_out_wire                 : std_logic_vector(31 downto 0); -- localedgepreserve_Fusion_Cal_Weight_0:max_out -> Bus_Conversion3:input
	signal localedgepreserve_fusion_cal_weight_0_value_out_wire               : std_logic_vector(31 downto 0); -- localedgepreserve_Fusion_Cal_Weight_0:value_out -> Bus_Conversion2:input
	signal localedgepreserve_fusion_cal_magnitude_gradient_2_0_valid_out_wire : std_logic;                     -- localedgepreserve_Fusion_Cal_Magnitude_Gradient_2_0:valid_out -> localedgepreserve_Fusion_Cal_A_B_2_0:valid_in
	signal valid1_in_0_output_wire                                            : std_logic;                     -- valid1_in_0:output -> localedgepreserve_Fusion_Cal_Magnitude_Gradient_1_0:valid_in
	signal pixel_in_0_output_wire                                             : std_logic_vector(7 downto 0);  -- pixel_in_0:output -> localedgepreserve_Fusion_Cal_Weight_0:pixel_in
	signal valid_in_0_output_wire                                             : std_logic;                     -- valid_in_0:output -> localedgepreserve_Fusion_Cal_Weight_0:valid_in
	signal eof_in_0_output_wire                                               : std_logic;                     -- eof_in_0:output -> localedgepreserve_Fusion_Cal_Weight_0:eof_in
	signal localedgepreserve_fusion_cal_image_out_2_0_ir_wire                 : std_logic_vector(7 downto 0);  -- localedgepreserve_Fusion_Cal_Image_Out_2_0:ir -> localedgepreserve_Fusion_Cal_Weight_0:addr_in
	signal eof1_in_0_output_wire                                              : std_logic;                     -- eof1_in_0:output -> localedgepreserve_Fusion_Cal_Magnitude_Gradient_1_0:eof_in
	signal localedgepreserve_fusion_cal_a_b_1_0_a_out_wire                    : std_logic_vector(15 downto 0); -- localedgepreserve_Fusion_Cal_A_B_1_0:a_out -> localedgepreserve_Fusion_Cal_Image_Out_1_0:a_in
	signal localedgepreserve_fusion_cal_a_b_1_0_valid_out_wire                : std_logic;                     -- localedgepreserve_Fusion_Cal_A_B_1_0:valid_out -> localedgepreserve_Fusion_Cal_Image_Out_1_0:valid_in
	signal localedgepreserve_fusion_cal_magnitude_gradient_1_0_valid_out_wire : std_logic;                     -- localedgepreserve_Fusion_Cal_Magnitude_Gradient_1_0:valid_out -> localedgepreserve_Fusion_Cal_A_B_1_0:valid_in
	signal localedgepreserve_fusion_cal_magnitude_gradient_1_0_eof_out_wire   : std_logic;                     -- localedgepreserve_Fusion_Cal_Magnitude_Gradient_1_0:eof_out -> localedgepreserve_Fusion_Cal_A_B_1_0:eof_in
	signal localedgepreserve_fusion_cal_a_b_1_0_b_out_wire                    : std_logic_vector(15 downto 0); -- localedgepreserve_Fusion_Cal_A_B_1_0:b_out -> localedgepreserve_Fusion_Cal_Image_Out_1_0:b_in
	signal localedgepreserve_fusion_cal_magnitude_gradient_2_0_eof_out_wire   : std_logic;                     -- localedgepreserve_Fusion_Cal_Magnitude_Gradient_2_0:eof_out -> localedgepreserve_Fusion_Cal_A_B_2_0:eof_in
	signal localedgepreserve_fusion_cal_a_b_2_0_b_out_wire                    : std_logic_vector(15 downto 0); -- localedgepreserve_Fusion_Cal_A_B_2_0:b_out -> localedgepreserve_Fusion_Cal_Image_Out_2_0:b_in
	signal localedgepreserve_fusion_cal_image_out_2_0_p_ir_wire               : std_logic_vector(15 downto 0); -- localedgepreserve_Fusion_Cal_Image_Out_2_0:p_ir -> Memory_Delay:input
	signal localedgepreserve_fusion_cal_image_out_1_0_p_vis_wire              : std_logic_vector(15 downto 0); -- localedgepreserve_Fusion_Cal_Image_Out_1_0:p_vis -> Memory_Delay1:input
	signal bus_conversion_output_wire                                         : std_logic_vector(8 downto 0);  -- Bus_Conversion:output -> [Multiplexer:in0, cast282:input]
	signal constant4_output_wire                                              : std_logic_vector(16 downto 0); -- Constant4:output -> Multiplexer1:in1
	signal memory_delay_output_wire                                           : std_logic_vector(15 downto 0); -- Memory_Delay:output -> Multiplier:datab
	signal multiplier_result_wire                                             : std_logic_vector(23 downto 0); -- Multiplier:result -> Delay:input
	signal multiplexer1_result_wire                                           : std_logic_vector(16 downto 0); -- Multiplexer1:result -> Multiplier1:dataa
	signal memory_delay1_output_wire                                          : std_logic_vector(15 downto 0); -- Memory_Delay1:output -> Multiplier1:datab
	signal constant_1_output_wire                                             : std_logic_vector(16 downto 0); -- Constant_1:output -> Pipelined_Adder:dataa
	signal pipelined_adder_result_wire                                        : std_logic_vector(16 downto 0); -- Pipelined_Adder:result -> Multiplexer1:in0
	signal pipelined_adder1_result_wire                                       : std_logic_vector(24 downto 0); -- Pipelined_Adder1:result -> Bus_Conversion:input
	signal localedgepreserve_fusion_cal_a_b_2_0_eof_out_wire                  : std_logic;                     -- localedgepreserve_Fusion_Cal_A_B_2_0:eof_out -> localedgepreserve_Fusion_generate_signals_0:eof_in
	signal multiplexer_result_wire                                            : std_logic_vector(8 downto 0);  -- Multiplexer:result -> pixel_out_0:input
	signal localedgepreserve_fusion_generate_signals_0_valid_out_wire         : std_logic;                     -- localedgepreserve_Fusion_generate_signals_0:valid_out -> valid_out_0:input
	signal localedgepreserve_fusion_generate_signals_0_sof_out_wire           : std_logic;                     -- localedgepreserve_Fusion_generate_signals_0:sof_out -> sof_out_0:input
	signal localedgepreserve_fusion_generate_signals_0_eof_out_wire           : std_logic;                     -- localedgepreserve_Fusion_generate_signals_0:eof_out -> eof_out_0:input
	signal binary_point_casting3_output_wire                                  : std_logic_vector(23 downto 0); -- Binary_Point_Casting3:output -> cast281:input
	signal cast281_output_wire                                                : std_logic_vector(23 downto 0); -- cast281:output -> Bus_Concatenation2:a
	signal cast282_output_wire                                                : std_logic_vector(9 downto 0);  -- cast282:output -> Comparator:dataa
	signal constant1_output_wire                                              : std_logic_vector(8 downto 0);  -- Constant1:output -> cast283:input
	signal cast283_output_wire                                                : std_logic_vector(9 downto 0);  -- cast283:output -> Comparator:datab
	signal constant3_output_wire                                              : std_logic_vector(16 downto 0); -- Constant3:output -> cast284:input
	signal cast284_output_wire                                                : std_logic_vector(17 downto 0); -- cast284:output -> Comparator1:datab
	signal delay1_output_wire                                                 : std_logic_vector(16 downto 0); -- Delay1:output -> cast285:input
	signal cast285_output_wire                                                : std_logic_vector(17 downto 0); -- cast285:output -> Comparator1:dataa
	signal bus_concatenation3_output_wire                                     : std_logic_vector(47 downto 0); -- Bus_Concatenation3:output -> cast286:input
	signal cast286_output_wire                                                : std_logic_vector(47 downto 0); -- cast286:output -> Divider:z
	signal binary_point_casting2_output_wire                                  : std_logic_vector(23 downto 0); -- Binary_Point_Casting2:output -> cast287:input
	signal cast287_output_wire                                                : std_logic_vector(23 downto 0); -- cast287:output -> Divider:d
	signal divider_q_wire                                                     : std_logic_vector(23 downto 0); -- Divider:q -> cast288:input
	signal cast288_output_wire                                                : std_logic_vector(23 downto 0); -- cast288:output -> Binary_Point_Casting1:input
	signal comparator_result_wire                                             : std_logic;                     -- Comparator:result -> cast289:input
	signal cast289_output_wire                                                : std_logic_vector(0 downto 0);  -- cast289:output -> Multiplexer:sel
	signal constant2_output_wire                                              : std_logic_vector(7 downto 0);  -- Constant2:output -> cast290:input
	signal cast290_output_wire                                                : std_logic_vector(8 downto 0);  -- cast290:output -> Multiplexer:in1
	signal comparator1_result_wire                                            : std_logic;                     -- Comparator1:result -> cast291:input
	signal cast291_output_wire                                                : std_logic_vector(0 downto 0);  -- cast291:output -> Multiplexer1:sel
	signal delay_output_wire                                                  : std_logic_vector(23 downto 0); -- Delay:output -> cast292:input
	signal cast292_output_wire                                                : std_logic_vector(24 downto 0); -- cast292:output -> Pipelined_Adder1:dataa
	signal multiplier1_result_wire                                            : std_logic_vector(23 downto 0); -- Multiplier1:result -> cast293:input
	signal cast293_output_wire                                                : std_logic_vector(24 downto 0); -- cast293:output -> Pipelined_Adder1:datab
	signal clock_0_clock_output_clk                                           : std_logic;                     -- Clock_0:clock_out -> [Bus_Concatenation2:clock, Bus_Concatenation3:clock, Comparator1:clock, Comparator:clock, Delay1:clock, Delay:clock, Divider:clk, Memory_Delay1:clock, Memory_Delay:clock, Multiplexer1:clock, Multiplexer:clock, Multiplier1:clock, Multiplier:clock, Pipelined_Adder1:clock, Pipelined_Adder:clock, localedgepreserve_Fusion_Cal_A_B_1_0:Clock, localedgepreserve_Fusion_Cal_A_B_2_0:Clock, localedgepreserve_Fusion_Cal_Image_Out_1_0:Clock, localedgepreserve_Fusion_Cal_Image_Out_2_0:Clock, localedgepreserve_Fusion_Cal_Magnitude_Gradient_1_0:Clock, localedgepreserve_Fusion_Cal_Magnitude_Gradient_2_0:Clock, localedgepreserve_Fusion_Cal_Weight_0:Clock, localedgepreserve_Fusion_generate_signals_0:Clock]
	signal clock_0_clock_output_reset                                         : std_logic;                     -- Clock_0:aclr_out -> [Bus_Concatenation2:aclr, Bus_Concatenation3:aclr, Comparator1:sclr, Comparator:sclr, Delay1:aclr, Delay:aclr, Memory_Delay1:aclr, Memory_Delay:aclr, Multiplexer1:aclr, Multiplexer:aclr, Multiplier1:aclr, Multiplier:aclr, Pipelined_Adder1:aclr, Pipelined_Adder:aclr, localedgepreserve_Fusion_Cal_A_B_1_0:reset, localedgepreserve_Fusion_Cal_A_B_2_0:reset, localedgepreserve_Fusion_Cal_Image_Out_1_0:reset, localedgepreserve_Fusion_Cal_Image_Out_2_0:reset, localedgepreserve_Fusion_Cal_Magnitude_Gradient_1_0:reset, localedgepreserve_Fusion_Cal_Magnitude_Gradient_2_0:reset, localedgepreserve_Fusion_Cal_Weight_0:reset, localedgepreserve_Fusion_generate_signals_0:reset]

begin

	clock_0 : component alt_dspbuilder_clock_GNQFU4PUDH
		port map (
			clock_out => clock_0_clock_output_clk,   -- clock_output.clk
			aclr_out  => clock_0_clock_output_reset, --             .reset
			clock     => Clock,                      --        clock.clk
			aclr      => reset                       --             .reset
		);

	valid_in_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => valid_in,               --  input.wire
			output => valid_in_0_output_wire  -- output.wire
		);

	multiplier1 : component alt_dspbuilder_multiplier_GNSFKO7633
		generic map (
			aWidth                         => 17,
			Signed                         => 0,
			bWidth                         => 16,
			DEDICATED_MULTIPLIER_CIRCUITRY => "YES",
			pipeline                       => 1,
			OutputLsb                      => 8,
			OutputMsb                      => 31
		)
		port map (
			clock     => clock_0_clock_output_clk,                            -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,                          --           .reset
			dataa     => multiplexer1_result_wire,                            --      dataa.wire
			datab     => memory_delay1_output_wire,                           --      datab.wire
			result    => multiplier1_result_wire,                             --     result.wire
			user_aclr => multiplier1user_aclrgnd_output_wire,                 --  user_aclr.wire
			ena       => localedgepreserve_fusion_cal_a_b_2_0_valid_out_wire  --        ena.wire
		);

	multiplier1user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplier1user_aclrgnd_output_wire  -- output.wire
		);

	binary_point_casting1 : component alt_dspbuilder_cast_GNUYRTQ4QH
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => cast288_output_wire,               --  input.wire
			output => binary_point_casting1_output_wire  -- output.wire
		);

	eof_out_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => localedgepreserve_fusion_generate_signals_0_eof_out_wire, --  input.wire
			output => eof_out                                                   -- output.wire
		);

	binary_point_casting3 : component alt_dspbuilder_cast_GNUYRTQ4QH
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => bus_conversion2_output_wire,       --  input.wire
			output => binary_point_casting3_output_wire  -- output.wire
		);

	binary_point_casting2 : component alt_dspbuilder_cast_GNUYRTQ4QH
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => bus_conversion3_output_wire,       --  input.wire
			output => binary_point_casting2_output_wire  -- output.wire
		);

	multiplexer : component alt_dspbuilder_multiplexer_GNIM5IEXF4
		generic map (
			number_inputs          => 2,
			pipeline               => 0,
			width                  => 9,
			HDLTYPE                => "STD_LOGIC_VECTOR",
			use_one_hot_select_bus => 0
		)
		port map (
			clock     => clock_0_clock_output_clk,            -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,          --           .reset
			sel       => cast289_output_wire,                 --        sel.wire
			result    => multiplexer_result_wire,             --     result.wire
			ena       => multiplexerenavcc_output_wire,       --        ena.wire
			user_aclr => multiplexeruser_aclrgnd_output_wire, --  user_aclr.wire
			in0       => bus_conversion_output_wire,          --        in0.wire
			in1       => cast290_output_wire                  --        in1.wire
		);

	multiplexeruser_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplexeruser_aclrgnd_output_wire  -- output.wire
		);

	multiplexerenavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => multiplexerenavcc_output_wire  -- output.wire
		);

	pixel_in_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => pixel_in,               --  input.wire
			output => pixel_in_0_output_wire  -- output.wire
		);

	localedgepreserve_fusion_cal_image_out_2_0 : component localedgepreserve_GN_localedgepreserve_Fusion_Cal_Image_Out_2
		port map (
			pixel_in => localedgepreserve_fusion_cal_a_b_2_0_pixel_out_wire,  -- pixel_in.wire
			a_in     => localedgepreserve_fusion_cal_a_b_2_0_a_out_wire,      --     a_in.wire
			b_in     => localedgepreserve_fusion_cal_a_b_2_0_b_out_wire,      --     b_in.wire
			ir       => localedgepreserve_fusion_cal_image_out_2_0_ir_wire,   --       ir.wire
			p_ir     => localedgepreserve_fusion_cal_image_out_2_0_p_ir_wire, --     p_ir.wire
			Clock    => clock_0_clock_output_clk,                             --    Clock.clk
			reset    => clock_0_clock_output_reset,                           --         .reset
			valid_in => localedgepreserve_fusion_cal_a_b_2_0_valid_out_wire   -- valid_in.wire
		);

	valid2_in_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => valid2_in,               --  input.wire
			output => valid2_in_0_output_wire  -- output.wire
		);

	delay : component alt_dspbuilder_delay_GNCY3KEQXH
		generic map (
			ClockPhase => "1",
			BitPattern => "000000010000000000000000",
			width      => 24,
			use_init   => 0,
			delay      => 1
		)
		port map (
			input  => multiplier_result_wire,                              --      input.wire
			clock  => clock_0_clock_output_clk,                            -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,                          --           .reset
			output => delay_output_wire,                                   --     output.wire
			sclr   => delaysclrgnd_output_wire,                            --       sclr.wire
			ena    => localedgepreserve_fusion_cal_a_b_2_0_valid_out_wire  --        ena.wire
		);

	delaysclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delaysclrgnd_output_wire  -- output.wire
		);

	localedgepreserve_fusion_cal_image_out_1_0 : component localedgepreserve_GN_localedgepreserve_Fusion_Cal_Image_Out_1
		port map (
			valid_in => localedgepreserve_fusion_cal_a_b_1_0_valid_out_wire,   -- valid_in.wire
			p_vis    => localedgepreserve_fusion_cal_image_out_1_0_p_vis_wire, --    p_vis.wire
			a_in     => localedgepreserve_fusion_cal_a_b_1_0_a_out_wire,       --     a_in.wire
			pixel_in => localedgepreserve_fusion_cal_a_b_1_0_pixel_out_wire,   -- pixel_in.wire
			Clock    => clock_0_clock_output_clk,                              --    Clock.clk
			reset    => clock_0_clock_output_reset,                            --         .reset
			b_in     => localedgepreserve_fusion_cal_a_b_1_0_b_out_wire        --     b_in.wire
		);

	comparator : component alt_dspbuilder_comparator_GN
		generic map (
			Operator  => "Altagb",
			lpm_width => 10
		)
		port map (
			clock  => clock_0_clock_output_clk,   -- clock_sclr.clk
			sclr   => clock_0_clock_output_reset, --           .reset
			dataa  => cast282_output_wire,        --      dataa.wire
			datab  => cast283_output_wire,        --      datab.wire
			result => comparator_result_wire      --     result.wire
		);

	localedgepreserve_fusion_generate_signals_0 : component localedgepreserve_GN_localedgepreserve_Fusion_generate_signals
		port map (
			eof_in    => localedgepreserve_fusion_cal_a_b_2_0_eof_out_wire,          --    eof_in.wire
			sof_out   => localedgepreserve_fusion_generate_signals_0_sof_out_wire,   --   sof_out.wire
			valid_in  => localedgepreserve_fusion_cal_a_b_2_0_valid_out_wire,        --  valid_in.wire
			valid_out => localedgepreserve_fusion_generate_signals_0_valid_out_wire, -- valid_out.wire
			Clock     => clock_0_clock_output_clk,                                   --     Clock.clk
			reset     => clock_0_clock_output_reset,                                 --          .reset
			eof_out   => localedgepreserve_fusion_generate_signals_0_eof_out_wire    --   eof_out.wire
		);

	eof1_in_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => eof1_in,               --  input.wire
			output => eof1_in_0_output_wire  -- output.wire
		);

	pipelined_adder1 : component alt_dspbuilder_pipelined_adder_GNTWZRTG4I
		generic map (
			pipeline => 1,
			width    => 25
		)
		port map (
			clock     => clock_0_clock_output_clk,                            -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,                          --           .reset
			dataa     => cast292_output_wire,                                 --      dataa.wire
			datab     => cast293_output_wire,                                 --      datab.wire
			result    => pipelined_adder1_result_wire,                        --     result.wire
			user_aclr => pipelined_adder1user_aclrgnd_output_wire,            --  user_aclr.wire
			ena       => localedgepreserve_fusion_cal_a_b_2_0_valid_out_wire  --        ena.wire
		);

	pipelined_adder1user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => pipelined_adder1user_aclrgnd_output_wire  -- output.wire
		);

	bus_conversion3 : component alt_dspbuilder_cast_GNEBWH7Z3U
		generic map (
			round    => 1,
			saturate => 0
		)
		port map (
			input  => localedgepreserve_fusion_cal_weight_0_max_out_wire, --  input.wire
			output => bus_conversion3_output_wire                         -- output.wire
		);

	bus_conversion2 : component alt_dspbuilder_cast_GNEBWH7Z3U
		generic map (
			round    => 1,
			saturate => 0
		)
		port map (
			input  => localedgepreserve_fusion_cal_weight_0_value_out_wire, --  input.wire
			output => bus_conversion2_output_wire                           -- output.wire
		);

	bus_conversion : component alt_dspbuilder_cast_GN7IYG3D6O
		generic map (
			round    => 1,
			saturate => 0
		)
		port map (
			input  => pipelined_adder1_result_wire, --  input.wire
			output => bus_conversion_output_wire    -- output.wire
		);

	bus_conversion1 : component alt_dspbuilder_cast_GNEL6FJM3V
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => binary_point_casting1_output_wire, --  input.wire
			output => bus_conversion1_output_wire        -- output.wire
		);

	constant2 : component alt_dspbuilder_constant_GNSVSRQZMI
		generic map (
			BitPattern => "11111111",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 8
		)
		port map (
			output => constant2_output_wire  -- output.wire
		);

	constant3 : component alt_dspbuilder_constant_GNQQLU6SNF
		generic map (
			BitPattern => "10000000000000000",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 17
		)
		port map (
			output => constant3_output_wire  -- output.wire
		);

	constant1 : component alt_dspbuilder_constant_GNP7U2HOAO
		generic map (
			BitPattern => "011111111",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 9
		)
		port map (
			output => constant1_output_wire  -- output.wire
		);

	valid1_in_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => valid1_in,               --  input.wire
			output => valid1_in_0_output_wire  -- output.wire
		);

	bus_concatenation2 : component alt_dspbuilder_bus_concat_GNU3KBQ5HN
		generic map (
			widthA => 24,
			widthB => 16
		)
		port map (
			clock  => clock_0_clock_output_clk,       -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,     --           .reset
			a      => cast281_output_wire,            --          a.wire
			b      => constant6_output_wire,          --          b.wire
			output => bus_concatenation2_output_wire  --     output.wire
		);

	bus_concatenation3 : component alt_dspbuilder_bus_concat_GN7K3OAUCY
		generic map (
			widthA => 8,
			widthB => 40
		)
		port map (
			clock  => clock_0_clock_output_clk,       -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,     --           .reset
			a      => constant7_output_wire,          --          a.wire
			b      => bus_concatenation2_output_wire, --          b.wire
			output => bus_concatenation3_output_wire  --     output.wire
		);

	constant6 : component alt_dspbuilder_constant_GNCWI5QDAD
		generic map (
			BitPattern => "0000000000000000",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 16
		)
		port map (
			output => constant6_output_wire  -- output.wire
		);

	constant7 : component alt_dspbuilder_constant_GNC5NOVIJT
		generic map (
			BitPattern => "00000000",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 8
		)
		port map (
			output => constant7_output_wire  -- output.wire
		);

	constant4 : component alt_dspbuilder_constant_GNDEA2MM7Q
		generic map (
			BitPattern => "00000000000000000",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 17
		)
		port map (
			output => constant4_output_wire  -- output.wire
		);

	sof_out_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => localedgepreserve_fusion_generate_signals_0_sof_out_wire, --  input.wire
			output => sof_out                                                   -- output.wire
		);

	eof2_in_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => eof2_in,               --  input.wire
			output => eof2_in_0_output_wire  -- output.wire
		);

	pixel_out_0 : component alt_dspbuilder_port_GNJVFJM3AT
		port map (
			input  => multiplexer_result_wire, --  input.wire
			output => pixel_out                -- output.wire
		);

	pixel2_in_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => pixel2_in,               --  input.wire
			output => pixel2_in_0_output_wire  -- output.wire
		);

	multiplexer1 : component alt_dspbuilder_multiplexer_GNMRY6PWYH
		generic map (
			number_inputs          => 2,
			pipeline               => 0,
			width                  => 17,
			HDLTYPE                => "STD_LOGIC_VECTOR",
			use_one_hot_select_bus => 0
		)
		port map (
			clock     => clock_0_clock_output_clk,             -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,           --           .reset
			sel       => cast291_output_wire,                  --        sel.wire
			result    => multiplexer1_result_wire,             --     result.wire
			ena       => multiplexer1enavcc_output_wire,       --        ena.wire
			user_aclr => multiplexer1user_aclrgnd_output_wire, --  user_aclr.wire
			in0       => pipelined_adder_result_wire,          --        in0.wire
			in1       => constant4_output_wire                 --        in1.wire
		);

	multiplexer1user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplexer1user_aclrgnd_output_wire  -- output.wire
		);

	multiplexer1enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => multiplexer1enavcc_output_wire  -- output.wire
		);

	localedgepreserve_fusion_cal_a_b_2_0 : component localedgepreserve_GN_localedgepreserve_Fusion_Cal_A_B_2
		port map (
			eof_in    => localedgepreserve_fusion_cal_magnitude_gradient_2_0_eof_out_wire,   --    eof_in.wire
			a_out     => localedgepreserve_fusion_cal_a_b_2_0_a_out_wire,                    --     a_out.wire
			pixel_in  => localedgepreserve_fusion_cal_magnitude_gradient_2_0_pixel_out_wire, --  pixel_in.wire
			b_out     => localedgepreserve_fusion_cal_a_b_2_0_b_out_wire,                    --     b_out.wire
			pixel_out => localedgepreserve_fusion_cal_a_b_2_0_pixel_out_wire,                -- pixel_out.wire
			Clock     => clock_0_clock_output_clk,                                           --     Clock.clk
			reset     => clock_0_clock_output_reset,                                         --          .reset
			grad_in   => localedgepreserve_fusion_cal_magnitude_gradient_2_0_grad_out_wire,  --   grad_in.wire
			eof_out   => localedgepreserve_fusion_cal_a_b_2_0_eof_out_wire,                  --   eof_out.wire
			valid_in  => localedgepreserve_fusion_cal_magnitude_gradient_2_0_valid_out_wire, --  valid_in.wire
			valid_out => localedgepreserve_fusion_cal_a_b_2_0_valid_out_wire                 -- valid_out.wire
		);

	pipelined_adder : component alt_dspbuilder_pipelined_adder_GNWEIMU3MK
		generic map (
			pipeline => 1,
			width    => 17
		)
		port map (
			clock     => clock_0_clock_output_clk,                            -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,                          --           .reset
			dataa     => constant_1_output_wire,                              --      dataa.wire
			datab     => bus_conversion1_output_wire,                         --      datab.wire
			result    => pipelined_adder_result_wire,                         --     result.wire
			user_aclr => pipelined_adderuser_aclrgnd_output_wire,             --  user_aclr.wire
			ena       => localedgepreserve_fusion_cal_a_b_2_0_valid_out_wire  --        ena.wire
		);

	pipelined_adderuser_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => pipelined_adderuser_aclrgnd_output_wire  -- output.wire
		);

	localedgepreserve_fusion_cal_a_b_1_0 : component localedgepreserve_GN_localedgepreserve_Fusion_Cal_A_B_1
		port map (
			eof_in    => localedgepreserve_fusion_cal_magnitude_gradient_1_0_eof_out_wire,   --    eof_in.wire
			b_out     => localedgepreserve_fusion_cal_a_b_1_0_b_out_wire,                    --     b_out.wire
			valid_out => localedgepreserve_fusion_cal_a_b_1_0_valid_out_wire,                -- valid_out.wire
			a_out     => localedgepreserve_fusion_cal_a_b_1_0_a_out_wire,                    --     a_out.wire
			pixel_out => localedgepreserve_fusion_cal_a_b_1_0_pixel_out_wire,                -- pixel_out.wire
			grad_in   => localedgepreserve_fusion_cal_magnitude_gradient_1_0_grad_out_wire,  --   grad_in.wire
			valid_in  => localedgepreserve_fusion_cal_magnitude_gradient_1_0_valid_out_wire, --  valid_in.wire
			pixel_in  => localedgepreserve_fusion_cal_magnitude_gradient_1_0_pixel_out_wire, --  pixel_in.wire
			Clock     => clock_0_clock_output_clk,                                           --     Clock.clk
			reset     => clock_0_clock_output_reset                                          --          .reset
		);

	comparator1 : component alt_dspbuilder_comparator_GN
		generic map (
			Operator  => "Altagb",
			lpm_width => 18
		)
		port map (
			clock  => clock_0_clock_output_clk,   -- clock_sclr.clk
			sclr   => clock_0_clock_output_reset, --           .reset
			dataa  => cast285_output_wire,        --      dataa.wire
			datab  => cast284_output_wire,        --      datab.wire
			result => comparator1_result_wire     --     result.wire
		);

	valid_out_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => localedgepreserve_fusion_generate_signals_0_valid_out_wire, --  input.wire
			output => valid_out                                                   -- output.wire
		);

	memory_delay1 : component alt_dspbuilder_memdelay_GNBRIKDQTV
		generic map (
			RAMTYPE => "AUTO",
			WIDTH   => 16,
			DELAY   => 26
		)
		port map (
			clock     => clock_0_clock_output_clk,                              -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,                            --           .reset
			input     => localedgepreserve_fusion_cal_image_out_1_0_p_vis_wire, --      input.wire
			output    => memory_delay1_output_wire,                             --     output.wire
			user_aclr => memory_delay1user_aclrgnd_output_wire,                 --  user_aclr.wire
			ena       => localedgepreserve_fusion_cal_a_b_2_0_valid_out_wire    --        ena.wire
		);

	memory_delay1user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => memory_delay1user_aclrgnd_output_wire  -- output.wire
		);

	multiplier : component alt_dspbuilder_multiplier_GNSFKO7633
		generic map (
			aWidth                         => 17,
			Signed                         => 0,
			bWidth                         => 16,
			DEDICATED_MULTIPLIER_CIRCUITRY => "YES",
			pipeline                       => 1,
			OutputLsb                      => 8,
			OutputMsb                      => 31
		)
		port map (
			clock     => clock_0_clock_output_clk,                            -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,                          --           .reset
			dataa     => bus_conversion1_output_wire,                         --      dataa.wire
			datab     => memory_delay_output_wire,                            --      datab.wire
			result    => multiplier_result_wire,                              --     result.wire
			user_aclr => multiplieruser_aclrgnd_output_wire,                  --  user_aclr.wire
			ena       => localedgepreserve_fusion_cal_a_b_2_0_valid_out_wire  --        ena.wire
		);

	multiplieruser_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplieruser_aclrgnd_output_wire  -- output.wire
		);

	pixel1_in_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => pixel1_in,               --  input.wire
			output => pixel1_in_0_output_wire  -- output.wire
		);

	delay1 : component alt_dspbuilder_delay_GNIDQK4WDH
		generic map (
			ClockPhase => "1",
			BitPattern => "10000000000000000",
			width      => 17,
			use_init   => 0,
			delay      => 1
		)
		port map (
			input  => bus_conversion1_output_wire,                         --      input.wire
			clock  => clock_0_clock_output_clk,                            -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,                          --           .reset
			output => delay1_output_wire,                                  --     output.wire
			sclr   => delay1sclrgnd_output_wire,                           --       sclr.wire
			ena    => localedgepreserve_fusion_cal_a_b_2_0_valid_out_wire  --        ena.wire
		);

	delay1sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delay1sclrgnd_output_wire  -- output.wire
		);

	localedgepreserve_fusion_cal_weight_0 : component localedgepreserve_GN_localedgepreserve_Fusion_Cal_Weight
		port map (
			max_out   => localedgepreserve_fusion_cal_weight_0_max_out_wire,   --   max_out.wire
			pixel_in  => pixel_in_0_output_wire,                               --  pixel_in.wire
			eof_in    => eof_in_0_output_wire,                                 --    eof_in.wire
			valid_in  => valid_in_0_output_wire,                               --  valid_in.wire
			value_out => localedgepreserve_fusion_cal_weight_0_value_out_wire, -- value_out.wire
			Clock     => clock_0_clock_output_clk,                             --     Clock.clk
			reset     => clock_0_clock_output_reset,                           --          .reset
			addr_in   => localedgepreserve_fusion_cal_image_out_2_0_ir_wire    --   addr_in.wire
		);

	eof_in_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => eof_in,               --  input.wire
			output => eof_in_0_output_wire  -- output.wire
		);

	localedgepreserve_fusion_cal_magnitude_gradient_2_0 : component localedgepreserve_GN_localedgepreserve_Fusion_Cal_Magnitude_Gradient_2
		port map (
			sof_out   => open,                                                               --   sof_out.wire
			pixel_out => localedgepreserve_fusion_cal_magnitude_gradient_2_0_pixel_out_wire, -- pixel_out.wire
			eof_out   => localedgepreserve_fusion_cal_magnitude_gradient_2_0_eof_out_wire,   --   eof_out.wire
			pixel_in  => pixel2_in_0_output_wire,                                            --  pixel_in.wire
			grad_out  => localedgepreserve_fusion_cal_magnitude_gradient_2_0_grad_out_wire,  --  grad_out.wire
			valid_out => localedgepreserve_fusion_cal_magnitude_gradient_2_0_valid_out_wire, -- valid_out.wire
			valid_in  => valid2_in_0_output_wire,                                            --  valid_in.wire
			Clock     => clock_0_clock_output_clk,                                           --     Clock.clk
			reset     => clock_0_clock_output_reset,                                         --          .reset
			eof_in    => eof2_in_0_output_wire                                               --    eof_in.wire
		);

	localedgepreserve_fusion_cal_magnitude_gradient_1_0 : component localedgepreserve_GN_localedgepreserve_Fusion_Cal_Magnitude_Gradient_1
		port map (
			eof_in    => eof1_in_0_output_wire,                                              --    eof_in.wire
			grad_out  => localedgepreserve_fusion_cal_magnitude_gradient_1_0_grad_out_wire,  --  grad_out.wire
			pixel_out => localedgepreserve_fusion_cal_magnitude_gradient_1_0_pixel_out_wire, -- pixel_out.wire
			valid_in  => valid1_in_0_output_wire,                                            --  valid_in.wire
			eof_out   => localedgepreserve_fusion_cal_magnitude_gradient_1_0_eof_out_wire,   --   eof_out.wire
			Clock     => clock_0_clock_output_clk,                                           --     Clock.clk
			reset     => clock_0_clock_output_reset,                                         --          .reset
			pixel_in  => pixel1_in_0_output_wire,                                            --  pixel_in.wire
			valid_out => localedgepreserve_fusion_cal_magnitude_gradient_1_0_valid_out_wire  -- valid_out.wire
		);

	constant_1 : component alt_dspbuilder_constant_GNQQLU6SNF
		generic map (
			BitPattern => "10000000000000000",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 17
		)
		port map (
			output => constant_1_output_wire  -- output.wire
		);

	memory_delay : component alt_dspbuilder_memdelay_GN3YPLAG7W
		generic map (
			RAMTYPE => "AUTO",
			WIDTH   => 16,
			DELAY   => 25
		)
		port map (
			clock     => clock_0_clock_output_clk,                             -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,                           --           .reset
			input     => localedgepreserve_fusion_cal_image_out_2_0_p_ir_wire, --      input.wire
			output    => memory_delay_output_wire,                             --     output.wire
			user_aclr => memory_delayuser_aclrgnd_output_wire,                 --  user_aclr.wire
			ena       => localedgepreserve_fusion_cal_a_b_2_0_valid_out_wire   --        ena.wire
		);

	memory_delayuser_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => memory_delayuser_aclrgnd_output_wire  -- output.wire
		);

	divider : component div
		port map (
			clk => clock_0_clock_output_clk,                            -- clk.clk
			ena => localedgepreserve_fusion_cal_a_b_2_0_valid_out_wire, -- ena.wire
			z   => cast286_output_wire,                                 --   z.wire
			d   => cast287_output_wire,                                 --   d.wire
			q   => divider_q_wire                                       --   q.wire
		);

	cast281 : component alt_dspbuilder_cast_GNA5TAMWCZ
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => binary_point_casting3_output_wire, --  input.wire
			output => cast281_output_wire                -- output.wire
		);

	cast282 : component alt_dspbuilder_cast_GNPFJ7B3O7
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => bus_conversion_output_wire, --  input.wire
			output => cast282_output_wire         -- output.wire
		);

	cast283 : component alt_dspbuilder_cast_GNPFJ7B3O7
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => constant1_output_wire, --  input.wire
			output => cast283_output_wire    -- output.wire
		);

	cast284 : component alt_dspbuilder_cast_GN7YNIFSF6
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => constant3_output_wire, --  input.wire
			output => cast284_output_wire    -- output.wire
		);

	cast285 : component alt_dspbuilder_cast_GN7YNIFSF6
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => delay1_output_wire,  --  input.wire
			output => cast285_output_wire  -- output.wire
		);

	cast286 : component alt_dspbuilder_cast_GNKD3JEUSD
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => bus_concatenation3_output_wire, --  input.wire
			output => cast286_output_wire             -- output.wire
		);

	cast287 : component alt_dspbuilder_cast_GN5P6ORZXA
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => binary_point_casting2_output_wire, --  input.wire
			output => cast287_output_wire                -- output.wire
		);

	cast288 : component alt_dspbuilder_cast_GNEIIG67TZ
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => divider_q_wire,      --  input.wire
			output => cast288_output_wire  -- output.wire
		);

	cast289 : component alt_dspbuilder_cast_GN46N4UJ5S
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => comparator_result_wire, --  input.wire
			output => cast289_output_wire     -- output.wire
		);

	cast290 : component alt_dspbuilder_cast_GNXDXNUGW4
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => constant2_output_wire, --  input.wire
			output => cast290_output_wire    -- output.wire
		);

	cast291 : component alt_dspbuilder_cast_GN46N4UJ5S
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => comparator1_result_wire, --  input.wire
			output => cast291_output_wire      -- output.wire
		);

	cast292 : component alt_dspbuilder_cast_GNJ6DWMNK6
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => delay_output_wire,   --  input.wire
			output => cast292_output_wire  -- output.wire
		);

	cast293 : component alt_dspbuilder_cast_GNJ6DWMNK6
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => multiplier1_result_wire, --  input.wire
			output => cast293_output_wire      -- output.wire
		);

end architecture rtl; -- of localedgepreserve_GN_localedgepreserve_Fusion
