-- gaussian_ip_GN_gaussian_ip_Fusion_Decomposition_3_multiplier_accumulator.vhd

-- Generated using ACDS version 17.1 590

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity gaussian_ip_GN_gaussian_ip_Fusion_Decomposition_3_multiplier_accumulator is
	port (
		pixel_out  : out std_logic_vector(31 downto 0);                    --  pixel_out.wire
		data_03    : in  std_logic_vector(7 downto 0)  := (others => '0'); --    data_03.wire
		data_43    : in  std_logic_vector(7 downto 0)  := (others => '0'); --    data_43.wire
		data_13    : in  std_logic_vector(7 downto 0)  := (others => '0'); --    data_13.wire
		data_30    : in  std_logic_vector(7 downto 0)  := (others => '0'); --    data_30.wire
		data_41    : in  std_logic_vector(7 downto 0)  := (others => '0'); --    data_41.wire
		clken      : in  std_logic                     := '0';             --      clken.wire
		data_12    : in  std_logic_vector(7 downto 0)  := (others => '0'); --    data_12.wire
		data_21    : in  std_logic_vector(7 downto 0)  := (others => '0'); --    data_21.wire
		Clock      : in  std_logic                     := '0';             --      Clock.clk
		reset      : in  std_logic                     := '0';             --           .reset
		data_23    : in  std_logic_vector(7 downto 0)  := (others => '0'); --    data_23.wire
		data_00    : in  std_logic_vector(7 downto 0)  := (others => '0'); --    data_00.wire
		data_11    : in  std_logic_vector(7 downto 0)  := (others => '0'); --    data_11.wire
		pixel_diff : out std_logic_vector(9 downto 0);                     -- pixel_diff.wire
		data_22    : in  std_logic_vector(7 downto 0)  := (others => '0'); --    data_22.wire
		data_24    : in  std_logic_vector(7 downto 0)  := (others => '0'); --    data_24.wire
		data_31    : in  std_logic_vector(7 downto 0)  := (others => '0'); --    data_31.wire
		data_02    : in  std_logic_vector(7 downto 0)  := (others => '0'); --    data_02.wire
		data_40    : in  std_logic_vector(7 downto 0)  := (others => '0'); --    data_40.wire
		data_33    : in  std_logic_vector(7 downto 0)  := (others => '0'); --    data_33.wire
		data_04    : in  std_logic_vector(7 downto 0)  := (others => '0'); --    data_04.wire
		data_32    : in  std_logic_vector(7 downto 0)  := (others => '0'); --    data_32.wire
		data_42    : in  std_logic_vector(7 downto 0)  := (others => '0'); --    data_42.wire
		data_10    : in  std_logic_vector(7 downto 0)  := (others => '0'); --    data_10.wire
		data_14    : in  std_logic_vector(7 downto 0)  := (others => '0'); --    data_14.wire
		data_20    : in  std_logic_vector(7 downto 0)  := (others => '0'); --    data_20.wire
		data_44    : in  std_logic_vector(7 downto 0)  := (others => '0'); --    data_44.wire
		data_34    : in  std_logic_vector(7 downto 0)  := (others => '0'); --    data_34.wire
		data_01    : in  std_logic_vector(7 downto 0)  := (others => '0')  --    data_01.wire
	);
end entity gaussian_ip_GN_gaussian_ip_Fusion_Decomposition_3_multiplier_accumulator;

architecture rtl of gaussian_ip_GN_gaussian_ip_Fusion_Decomposition_3_multiplier_accumulator is
	component alt_dspbuilder_clock_GNQFU4PUDH is
		port (
			aclr      : in  std_logic := 'X'; -- reset
			aclr_n    : in  std_logic := 'X'; -- reset_n
			aclr_out  : out std_logic;        -- reset
			clock     : in  std_logic := 'X'; -- clk
			clock_out : out std_logic         -- clk
		);
	end component alt_dspbuilder_clock_GNQFU4PUDH;

	component alt_dspbuilder_multiplier_GNNIEJHQ5V is
		generic (
			aWidth                         : natural := 8;
			Signed                         : natural := 0;
			bWidth                         : natural := 8;
			DEDICATED_MULTIPLIER_CIRCUITRY : string  := "AUTO";
			pipeline                       : integer := 0;
			OutputLsb                      : integer := 0;
			OutputMsb                      : integer := 8
		);
		port (
			aclr      : in  std_logic                                          := 'X';             -- clk
			clock     : in  std_logic                                          := 'X';             -- clk
			dataa     : in  std_logic_vector(aWidth-1 downto 0)                := (others => 'X'); -- wire
			datab     : in  std_logic_vector(bWidth-1 downto 0)                := (others => 'X'); -- wire
			ena       : in  std_logic                                          := 'X';             -- wire
			result    : out std_logic_vector(OutputMsb-OutputLsb+1-1 downto 0);                    -- wire
			user_aclr : in  std_logic                                          := 'X'              -- wire
		);
	end component alt_dspbuilder_multiplier_GNNIEJHQ5V;

	component alt_dspbuilder_gnd_GN is
		port (
			output : out std_logic   -- wire
		);
	end component alt_dspbuilder_gnd_GN;

	component alt_dspbuilder_constant_GN6SFEINY6 is
		generic (
			BitPattern : string  := "0000";
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(1 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GN6SFEINY6;

	component alt_dspbuilder_constant_GN2DUUMQHA is
		generic (
			BitPattern : string  := "0000";
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(25 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GN2DUUMQHA;

	component alt_dspbuilder_constant_GN52UV6F2X is
		generic (
			BitPattern : string  := "0000";
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(25 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GN52UV6F2X;

	component alt_dspbuilder_constant_GNBQQQV5ZM is
		generic (
			BitPattern : string  := "0000";
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(25 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GNBQQQV5ZM;

	component alt_dspbuilder_port_GNA5S4SQDN is
		port (
			input  : in  std_logic_vector(7 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(7 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNA5S4SQDN;

	component alt_dspbuilder_bus_concat_GNKLOJ6ING is
		generic (
			widthA : natural := 8;
			widthB : natural := 8
		);
		port (
			a      : in  std_logic_vector(widthA-1 downto 0)        := (others => 'X'); -- wire
			aclr   : in  std_logic                                  := 'X';             -- clk
			b      : in  std_logic_vector(widthB-1 downto 0)        := (others => 'X'); -- wire
			clock  : in  std_logic                                  := 'X';             -- clk
			output : out std_logic_vector(widthA+widthB-1 downto 0)                     -- wire
		);
	end component alt_dspbuilder_bus_concat_GNKLOJ6ING;

	component alt_dspbuilder_constant_GN42V6LR6J is
		generic (
			BitPattern : string  := "0000";
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(25 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GN42V6LR6J;

	component alt_dspbuilder_constant_GN3UR3AYSK is
		generic (
			BitPattern : string  := "0000";
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(25 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GN3UR3AYSK;

	component alt_dspbuilder_port_GNEPKLLZKY is
		port (
			input  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(31 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNEPKLLZKY;

	component alt_dspbuilder_pipelined_adder_GNY2JEH574 is
		generic (
			pipeline : integer := 0;
			width    : natural := 0
		);
		port (
			aclr      : in  std_logic                          := 'X';             -- clk
			add_sub   : in  std_logic                          := 'X';             -- wire
			cin       : in  std_logic                          := 'X';             -- wire
			clock     : in  std_logic                          := 'X';             -- clk
			cout      : out std_logic;                                             -- wire
			dataa     : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			datab     : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			ena       : in  std_logic                          := 'X';             -- wire
			result    : out std_logic_vector(width-1 downto 0);                    -- wire
			user_aclr : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_pipelined_adder_GNY2JEH574;

	component alt_dspbuilder_port_GNSSYS4J5R is
		port (
			input  : in  std_logic_vector(9 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(9 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNSSYS4J5R;

	component alt_dspbuilder_round_GNWBUVGWWO is
		generic (
			OUT_WIDTH_g     : natural := 6;
			IN_WIDTH_g      : natural := 8;
			PIPELINE_g      : natural := 0;
			ROUNDING_TYPE_g : string  := "TRUNCATE_LOW";
			SIGNED_g        : natural := 1
		);
		port (
			clk       : in  std_logic                     := 'X';             -- clk
			reset     : in  std_logic                     := 'X';             -- wire
			datain    : in  std_logic_vector(25 downto 0) := (others => 'X'); -- wire
			dataout   : out std_logic_vector(7 downto 0);                     -- wire
			ena       : in  std_logic                     := 'X';             -- wire
			user_aclr : in  std_logic                     := 'X'              -- wire
		);
	end component alt_dspbuilder_round_GNWBUVGWWO;

	component alt_dspbuilder_vcc_GN is
		port (
			output : out std_logic   -- wire
		);
	end component alt_dspbuilder_vcc_GN;

	component alt_dspbuilder_parallel_adder_GN5CSCONM5 is
		generic (
			dataWidth     : positive := 8;
			direction     : string   := "+";
			MaskValue     : string   := "1";
			pipeline      : natural  := 0;
			number_inputs : positive := 2
		);
		port (
			clock     : in  std_logic                     := 'X';             -- clk
			aclr      : in  std_logic                     := 'X';             -- reset
			result    : out std_logic_vector(31 downto 0);                    -- wire
			user_aclr : in  std_logic                     := 'X';             -- wire
			ena       : in  std_logic                     := 'X';             -- wire
			data0     : in  std_logic_vector(26 downto 0) := (others => 'X'); -- wire
			data1     : in  std_logic_vector(26 downto 0) := (others => 'X'); -- wire
			data2     : in  std_logic_vector(26 downto 0) := (others => 'X'); -- wire
			data3     : in  std_logic_vector(26 downto 0) := (others => 'X'); -- wire
			data4     : in  std_logic_vector(26 downto 0) := (others => 'X'); -- wire
			data5     : in  std_logic_vector(26 downto 0) := (others => 'X'); -- wire
			data6     : in  std_logic_vector(26 downto 0) := (others => 'X'); -- wire
			data7     : in  std_logic_vector(26 downto 0) := (others => 'X'); -- wire
			data8     : in  std_logic_vector(26 downto 0) := (others => 'X'); -- wire
			data9     : in  std_logic_vector(26 downto 0) := (others => 'X'); -- wire
			data10    : in  std_logic_vector(26 downto 0) := (others => 'X'); -- wire
			data11    : in  std_logic_vector(26 downto 0) := (others => 'X'); -- wire
			data12    : in  std_logic_vector(26 downto 0) := (others => 'X'); -- wire
			data13    : in  std_logic_vector(26 downto 0) := (others => 'X'); -- wire
			data14    : in  std_logic_vector(26 downto 0) := (others => 'X'); -- wire
			data15    : in  std_logic_vector(26 downto 0) := (others => 'X'); -- wire
			data16    : in  std_logic_vector(26 downto 0) := (others => 'X'); -- wire
			data17    : in  std_logic_vector(26 downto 0) := (others => 'X'); -- wire
			data18    : in  std_logic_vector(26 downto 0) := (others => 'X'); -- wire
			data19    : in  std_logic_vector(26 downto 0) := (others => 'X'); -- wire
			data20    : in  std_logic_vector(26 downto 0) := (others => 'X'); -- wire
			data21    : in  std_logic_vector(26 downto 0) := (others => 'X'); -- wire
			data22    : in  std_logic_vector(26 downto 0) := (others => 'X'); -- wire
			data23    : in  std_logic_vector(26 downto 0) := (others => 'X'); -- wire
			data24    : in  std_logic_vector(26 downto 0) := (others => 'X')  -- wire
		);
	end component alt_dspbuilder_parallel_adder_GN5CSCONM5;

	component alt_dspbuilder_constant_GNHUGKQYBA is
		generic (
			BitPattern : string  := "0000";
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(25 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GNHUGKQYBA;

	component alt_dspbuilder_port_GN37ALZBS4 is
		port (
			input  : in  std_logic := 'X'; -- wire
			output : out std_logic         -- wire
		);
	end component alt_dspbuilder_port_GN37ALZBS4;

	component alt_dspbuilder_memdelay_GND4ZY57YF is
		generic (
			RAMTYPE : string   := "AUTO";
			WIDTH   : positive := 8;
			DELAY   : positive := 1
		);
		port (
			aclr      : in  std_logic                          := 'X';             -- clk
			clock     : in  std_logic                          := 'X';             -- clk
			ena       : in  std_logic                          := 'X';             -- wire
			input     : in  std_logic_vector(WIDTH-1 downto 0) := (others => 'X'); -- wire
			output    : out std_logic_vector(WIDTH-1 downto 0);                    -- wire
			user_aclr : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_memdelay_GND4ZY57YF;

	component alt_dspbuilder_cast_GNBZR5PMEK is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(7 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(7 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNBZR5PMEK;

	component alt_dspbuilder_cast_GNMLNX2RCD is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(25 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(26 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNMLNX2RCD;

	component alt_dspbuilder_cast_GNHYNEPC7U is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(25 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNHYNEPC7U;

	signal multiplier2user_aclrgnd_output_wire               : std_logic;                     -- Multiplier2user_aclrGND:output -> Multiplier2:user_aclr
	signal multiplier1user_aclrgnd_output_wire               : std_logic;                     -- Multiplier1user_aclrGND:output -> Multiplier1:user_aclr
	signal multiplier18user_aclrgnd_output_wire              : std_logic;                     -- Multiplier18user_aclrGND:output -> Multiplier18:user_aclr
	signal multiplier4user_aclrgnd_output_wire               : std_logic;                     -- Multiplier4user_aclrGND:output -> Multiplier4:user_aclr
	signal multiplier19user_aclrgnd_output_wire              : std_logic;                     -- Multiplier19user_aclrGND:output -> Multiplier19:user_aclr
	signal multiplier3user_aclrgnd_output_wire               : std_logic;                     -- Multiplier3user_aclrGND:output -> Multiplier3:user_aclr
	signal multiplier6user_aclrgnd_output_wire               : std_logic;                     -- Multiplier6user_aclrGND:output -> Multiplier6:user_aclr
	signal multiplier5user_aclrgnd_output_wire               : std_logic;                     -- Multiplier5user_aclrGND:output -> Multiplier5:user_aclr
	signal multiplier8user_aclrgnd_output_wire               : std_logic;                     -- Multiplier8user_aclrGND:output -> Multiplier8:user_aclr
	signal multiplier7user_aclrgnd_output_wire               : std_logic;                     -- Multiplier7user_aclrGND:output -> Multiplier7:user_aclr
	signal multiplier12user_aclrgnd_output_wire              : std_logic;                     -- Multiplier12user_aclrGND:output -> Multiplier12:user_aclr
	signal multiplier13user_aclrgnd_output_wire              : std_logic;                     -- Multiplier13user_aclrGND:output -> Multiplier13:user_aclr
	signal multiplier9user_aclrgnd_output_wire               : std_logic;                     -- Multiplier9user_aclrGND:output -> Multiplier9:user_aclr
	signal multiplier10user_aclrgnd_output_wire              : std_logic;                     -- Multiplier10user_aclrGND:output -> Multiplier10:user_aclr
	signal multiplier11user_aclrgnd_output_wire              : std_logic;                     -- Multiplier11user_aclrGND:output -> Multiplier11:user_aclr
	signal multiplier16user_aclrgnd_output_wire              : std_logic;                     -- Multiplier16user_aclrGND:output -> Multiplier16:user_aclr
	signal multiplier17user_aclrgnd_output_wire              : std_logic;                     -- Multiplier17user_aclrGND:output -> Multiplier17:user_aclr
	signal multiplier14user_aclrgnd_output_wire              : std_logic;                     -- Multiplier14user_aclrGND:output -> Multiplier14:user_aclr
	signal multiplier15user_aclrgnd_output_wire              : std_logic;                     -- Multiplier15user_aclrGND:output -> Multiplier15:user_aclr
	signal multiplier20user_aclrgnd_output_wire              : std_logic;                     -- Multiplier20user_aclrGND:output -> Multiplier20:user_aclr
	signal multiplier23user_aclrgnd_output_wire              : std_logic;                     -- Multiplier23user_aclrGND:output -> Multiplier23:user_aclr
	signal multiplier24user_aclrgnd_output_wire              : std_logic;                     -- Multiplier24user_aclrGND:output -> Multiplier24:user_aclr
	signal multiplier21user_aclrgnd_output_wire              : std_logic;                     -- Multiplier21user_aclrGND:output -> Multiplier21:user_aclr
	signal multiplier22user_aclrgnd_output_wire              : std_logic;                     -- Multiplier22user_aclrGND:output -> Multiplier22:user_aclr
	signal pipelined_adderuser_aclrgnd_output_wire           : std_logic;                     -- Pipelined_Adderuser_aclrGND:output -> Pipelined_Adder:user_aclr
	signal multiplieruser_aclrgnd_output_wire                : std_logic;                     -- Multiplieruser_aclrGND:output -> Multiplier:user_aclr
	signal rounduser_aclrgnd_output_wire                     : std_logic;                     -- Rounduser_aclrGND:output -> Round:user_aclr
	signal roundenavcc_output_wire                           : std_logic;                     -- RoundenaVCC:output -> Round:ena
	signal roundresetgnd_output_wire                         : std_logic;                     -- RoundresetGND:output -> Round:reset
	signal parallel_adder_subtractoruser_aclrgnd_output_wire : std_logic;                     -- Parallel_Adder_Subtractoruser_aclrGND:output -> Parallel_Adder_Subtractor:user_aclr
	signal memory_delayuser_aclrgnd_output_wire              : std_logic;                     -- Memory_Delayuser_aclrGND:output -> Memory_Delay:user_aclr
	signal constant25_output_wire                            : std_logic_vector(1 downto 0);  -- Constant25:output -> Bus_Concatenation1:a
	signal constant26_output_wire                            : std_logic_vector(1 downto 0);  -- Constant26:output -> Bus_Concatenation:a
	signal data_22_0_output_wire                             : std_logic_vector(7 downto 0);  -- data_22_0:output -> [Memory_Delay:input, Multiplier12:dataa]
	signal clken_0_output_wire                               : std_logic;                     -- clken_0:output -> [Memory_Delay:ena, Multiplier10:ena, Multiplier11:ena, Multiplier12:ena, Multiplier13:ena, Multiplier14:ena, Multiplier15:ena, Multiplier16:ena, Multiplier17:ena, Multiplier18:ena, Multiplier19:ena, Multiplier1:ena, Multiplier20:ena, Multiplier21:ena, Multiplier22:ena, Multiplier23:ena, Multiplier24:ena, Multiplier2:ena, Multiplier3:ena, Multiplier4:ena, Multiplier5:ena, Multiplier6:ena, Multiplier7:ena, Multiplier8:ena, Multiplier9:ena, Multiplier:ena, Parallel_Adder_Subtractor:ena, Pipelined_Adder:ena]
	signal data_00_0_output_wire                             : std_logic_vector(7 downto 0);  -- data_00_0:output -> Multiplier:dataa
	signal constant_1_output_wire                            : std_logic_vector(25 downto 0); -- Constant_1:output -> Multiplier:datab
	signal data_01_0_output_wire                             : std_logic_vector(7 downto 0);  -- data_01_0:output -> Multiplier1:dataa
	signal constant1_output_wire                             : std_logic_vector(25 downto 0); -- Constant1:output -> Multiplier1:datab
	signal data_20_0_output_wire                             : std_logic_vector(7 downto 0);  -- data_20_0:output -> Multiplier10:dataa
	signal constant10_output_wire                            : std_logic_vector(25 downto 0); -- Constant10:output -> Multiplier10:datab
	signal data_21_0_output_wire                             : std_logic_vector(7 downto 0);  -- data_21_0:output -> Multiplier11:dataa
	signal constant11_output_wire                            : std_logic_vector(25 downto 0); -- Constant11:output -> Multiplier11:datab
	signal constant12_output_wire                            : std_logic_vector(25 downto 0); -- Constant12:output -> Multiplier12:datab
	signal data_23_0_output_wire                             : std_logic_vector(7 downto 0);  -- data_23_0:output -> Multiplier13:dataa
	signal constant13_output_wire                            : std_logic_vector(25 downto 0); -- Constant13:output -> Multiplier13:datab
	signal data_24_0_output_wire                             : std_logic_vector(7 downto 0);  -- data_24_0:output -> Multiplier14:dataa
	signal constant14_output_wire                            : std_logic_vector(25 downto 0); -- Constant14:output -> Multiplier14:datab
	signal data_30_0_output_wire                             : std_logic_vector(7 downto 0);  -- data_30_0:output -> Multiplier15:dataa
	signal constant15_output_wire                            : std_logic_vector(25 downto 0); -- Constant15:output -> Multiplier15:datab
	signal data_31_0_output_wire                             : std_logic_vector(7 downto 0);  -- data_31_0:output -> Multiplier16:dataa
	signal constant16_output_wire                            : std_logic_vector(25 downto 0); -- Constant16:output -> Multiplier16:datab
	signal data_32_0_output_wire                             : std_logic_vector(7 downto 0);  -- data_32_0:output -> Multiplier17:dataa
	signal constant17_output_wire                            : std_logic_vector(25 downto 0); -- Constant17:output -> Multiplier17:datab
	signal data_33_0_output_wire                             : std_logic_vector(7 downto 0);  -- data_33_0:output -> Multiplier18:dataa
	signal constant18_output_wire                            : std_logic_vector(25 downto 0); -- Constant18:output -> Multiplier18:datab
	signal data_34_0_output_wire                             : std_logic_vector(7 downto 0);  -- data_34_0:output -> Multiplier19:dataa
	signal constant19_output_wire                            : std_logic_vector(25 downto 0); -- Constant19:output -> Multiplier19:datab
	signal data_02_0_output_wire                             : std_logic_vector(7 downto 0);  -- data_02_0:output -> Multiplier2:dataa
	signal constant2_output_wire                             : std_logic_vector(25 downto 0); -- Constant2:output -> Multiplier2:datab
	signal data_40_0_output_wire                             : std_logic_vector(7 downto 0);  -- data_40_0:output -> Multiplier20:dataa
	signal constant20_output_wire                            : std_logic_vector(25 downto 0); -- Constant20:output -> Multiplier20:datab
	signal data_41_0_output_wire                             : std_logic_vector(7 downto 0);  -- data_41_0:output -> Multiplier21:dataa
	signal constant21_output_wire                            : std_logic_vector(25 downto 0); -- Constant21:output -> Multiplier21:datab
	signal data_42_0_output_wire                             : std_logic_vector(7 downto 0);  -- data_42_0:output -> Multiplier22:dataa
	signal constant22_output_wire                            : std_logic_vector(25 downto 0); -- Constant22:output -> Multiplier22:datab
	signal data_43_0_output_wire                             : std_logic_vector(7 downto 0);  -- data_43_0:output -> Multiplier23:dataa
	signal constant23_output_wire                            : std_logic_vector(25 downto 0); -- Constant23:output -> Multiplier23:datab
	signal data_44_0_output_wire                             : std_logic_vector(7 downto 0);  -- data_44_0:output -> Multiplier24:dataa
	signal constant24_output_wire                            : std_logic_vector(25 downto 0); -- Constant24:output -> Multiplier24:datab
	signal data_03_0_output_wire                             : std_logic_vector(7 downto 0);  -- data_03_0:output -> Multiplier3:dataa
	signal constant3_output_wire                             : std_logic_vector(25 downto 0); -- Constant3:output -> Multiplier3:datab
	signal data_04_0_output_wire                             : std_logic_vector(7 downto 0);  -- data_04_0:output -> Multiplier4:dataa
	signal constant4_output_wire                             : std_logic_vector(25 downto 0); -- Constant4:output -> Multiplier4:datab
	signal data_10_0_output_wire                             : std_logic_vector(7 downto 0);  -- data_10_0:output -> Multiplier5:dataa
	signal constant5_output_wire                             : std_logic_vector(25 downto 0); -- Constant5:output -> Multiplier5:datab
	signal data_11_0_output_wire                             : std_logic_vector(7 downto 0);  -- data_11_0:output -> Multiplier6:dataa
	signal constant6_output_wire                             : std_logic_vector(25 downto 0); -- Constant6:output -> Multiplier6:datab
	signal data_12_0_output_wire                             : std_logic_vector(7 downto 0);  -- data_12_0:output -> Multiplier7:dataa
	signal constant7_output_wire                             : std_logic_vector(25 downto 0); -- Constant7:output -> Multiplier7:datab
	signal data_13_0_output_wire                             : std_logic_vector(7 downto 0);  -- data_13_0:output -> Multiplier8:dataa
	signal constant8_output_wire                             : std_logic_vector(25 downto 0); -- Constant8:output -> Multiplier8:datab
	signal data_14_0_output_wire                             : std_logic_vector(7 downto 0);  -- data_14_0:output -> Multiplier9:dataa
	signal constant9_output_wire                             : std_logic_vector(25 downto 0); -- Constant9:output -> Multiplier9:datab
	signal bus_concatenation1_output_wire                    : std_logic_vector(9 downto 0);  -- Bus_Concatenation1:output -> Pipelined_Adder:dataa
	signal bus_concatenation_output_wire                     : std_logic_vector(9 downto 0);  -- Bus_Concatenation:output -> Pipelined_Adder:datab
	signal parallel_adder_subtractor_result_wire             : std_logic_vector(31 downto 0); -- Parallel_Adder_Subtractor:result -> [cast26:input, pixel_out_0:input]
	signal pipelined_adder_result_wire                       : std_logic_vector(9 downto 0);  -- Pipelined_Adder:result -> pixel_diff_0:input
	signal memory_delay_output_wire                          : std_logic_vector(7 downto 0);  -- Memory_Delay:output -> cast0:input
	signal cast0_output_wire                                 : std_logic_vector(7 downto 0);  -- cast0:output -> Bus_Concatenation1:b
	signal multiplier_result_wire                            : std_logic_vector(25 downto 0); -- Multiplier:result -> cast1:input
	signal cast1_output_wire                                 : std_logic_vector(26 downto 0); -- cast1:output -> Parallel_Adder_Subtractor:data0
	signal multiplier1_result_wire                           : std_logic_vector(25 downto 0); -- Multiplier1:result -> cast2:input
	signal cast2_output_wire                                 : std_logic_vector(26 downto 0); -- cast2:output -> Parallel_Adder_Subtractor:data1
	signal multiplier2_result_wire                           : std_logic_vector(25 downto 0); -- Multiplier2:result -> cast3:input
	signal cast3_output_wire                                 : std_logic_vector(26 downto 0); -- cast3:output -> Parallel_Adder_Subtractor:data2
	signal multiplier3_result_wire                           : std_logic_vector(25 downto 0); -- Multiplier3:result -> cast4:input
	signal cast4_output_wire                                 : std_logic_vector(26 downto 0); -- cast4:output -> Parallel_Adder_Subtractor:data3
	signal multiplier4_result_wire                           : std_logic_vector(25 downto 0); -- Multiplier4:result -> cast5:input
	signal cast5_output_wire                                 : std_logic_vector(26 downto 0); -- cast5:output -> Parallel_Adder_Subtractor:data4
	signal multiplier5_result_wire                           : std_logic_vector(25 downto 0); -- Multiplier5:result -> cast6:input
	signal cast6_output_wire                                 : std_logic_vector(26 downto 0); -- cast6:output -> Parallel_Adder_Subtractor:data5
	signal multiplier6_result_wire                           : std_logic_vector(25 downto 0); -- Multiplier6:result -> cast7:input
	signal cast7_output_wire                                 : std_logic_vector(26 downto 0); -- cast7:output -> Parallel_Adder_Subtractor:data6
	signal multiplier7_result_wire                           : std_logic_vector(25 downto 0); -- Multiplier7:result -> cast8:input
	signal cast8_output_wire                                 : std_logic_vector(26 downto 0); -- cast8:output -> Parallel_Adder_Subtractor:data7
	signal multiplier8_result_wire                           : std_logic_vector(25 downto 0); -- Multiplier8:result -> cast9:input
	signal cast9_output_wire                                 : std_logic_vector(26 downto 0); -- cast9:output -> Parallel_Adder_Subtractor:data8
	signal multiplier9_result_wire                           : std_logic_vector(25 downto 0); -- Multiplier9:result -> cast10:input
	signal cast10_output_wire                                : std_logic_vector(26 downto 0); -- cast10:output -> Parallel_Adder_Subtractor:data9
	signal multiplier10_result_wire                          : std_logic_vector(25 downto 0); -- Multiplier10:result -> cast11:input
	signal cast11_output_wire                                : std_logic_vector(26 downto 0); -- cast11:output -> Parallel_Adder_Subtractor:data10
	signal multiplier11_result_wire                          : std_logic_vector(25 downto 0); -- Multiplier11:result -> cast12:input
	signal cast12_output_wire                                : std_logic_vector(26 downto 0); -- cast12:output -> Parallel_Adder_Subtractor:data11
	signal multiplier12_result_wire                          : std_logic_vector(25 downto 0); -- Multiplier12:result -> cast13:input
	signal cast13_output_wire                                : std_logic_vector(26 downto 0); -- cast13:output -> Parallel_Adder_Subtractor:data12
	signal multiplier13_result_wire                          : std_logic_vector(25 downto 0); -- Multiplier13:result -> cast14:input
	signal cast14_output_wire                                : std_logic_vector(26 downto 0); -- cast14:output -> Parallel_Adder_Subtractor:data13
	signal multiplier14_result_wire                          : std_logic_vector(25 downto 0); -- Multiplier14:result -> cast15:input
	signal cast15_output_wire                                : std_logic_vector(26 downto 0); -- cast15:output -> Parallel_Adder_Subtractor:data14
	signal multiplier15_result_wire                          : std_logic_vector(25 downto 0); -- Multiplier15:result -> cast16:input
	signal cast16_output_wire                                : std_logic_vector(26 downto 0); -- cast16:output -> Parallel_Adder_Subtractor:data15
	signal multiplier16_result_wire                          : std_logic_vector(25 downto 0); -- Multiplier16:result -> cast17:input
	signal cast17_output_wire                                : std_logic_vector(26 downto 0); -- cast17:output -> Parallel_Adder_Subtractor:data16
	signal multiplier17_result_wire                          : std_logic_vector(25 downto 0); -- Multiplier17:result -> cast18:input
	signal cast18_output_wire                                : std_logic_vector(26 downto 0); -- cast18:output -> Parallel_Adder_Subtractor:data17
	signal multiplier18_result_wire                          : std_logic_vector(25 downto 0); -- Multiplier18:result -> cast19:input
	signal cast19_output_wire                                : std_logic_vector(26 downto 0); -- cast19:output -> Parallel_Adder_Subtractor:data18
	signal multiplier19_result_wire                          : std_logic_vector(25 downto 0); -- Multiplier19:result -> cast20:input
	signal cast20_output_wire                                : std_logic_vector(26 downto 0); -- cast20:output -> Parallel_Adder_Subtractor:data19
	signal multiplier20_result_wire                          : std_logic_vector(25 downto 0); -- Multiplier20:result -> cast21:input
	signal cast21_output_wire                                : std_logic_vector(26 downto 0); -- cast21:output -> Parallel_Adder_Subtractor:data20
	signal multiplier21_result_wire                          : std_logic_vector(25 downto 0); -- Multiplier21:result -> cast22:input
	signal cast22_output_wire                                : std_logic_vector(26 downto 0); -- cast22:output -> Parallel_Adder_Subtractor:data21
	signal multiplier22_result_wire                          : std_logic_vector(25 downto 0); -- Multiplier22:result -> cast23:input
	signal cast23_output_wire                                : std_logic_vector(26 downto 0); -- cast23:output -> Parallel_Adder_Subtractor:data22
	signal multiplier23_result_wire                          : std_logic_vector(25 downto 0); -- Multiplier23:result -> cast24:input
	signal cast24_output_wire                                : std_logic_vector(26 downto 0); -- cast24:output -> Parallel_Adder_Subtractor:data23
	signal multiplier24_result_wire                          : std_logic_vector(25 downto 0); -- Multiplier24:result -> cast25:input
	signal cast25_output_wire                                : std_logic_vector(26 downto 0); -- cast25:output -> Parallel_Adder_Subtractor:data24
	signal cast26_output_wire                                : std_logic_vector(25 downto 0); -- cast26:output -> Round:datain
	signal round_dataout_wire                                : std_logic_vector(7 downto 0);  -- Round:dataout -> cast27:input
	signal cast27_output_wire                                : std_logic_vector(7 downto 0);  -- cast27:output -> Bus_Concatenation:b
	signal clock_0_clock_output_clk                          : std_logic;                     -- Clock_0:clock_out -> [Bus_Concatenation1:clock, Bus_Concatenation:clock, Memory_Delay:clock, Multiplier10:clock, Multiplier11:clock, Multiplier12:clock, Multiplier13:clock, Multiplier14:clock, Multiplier15:clock, Multiplier16:clock, Multiplier17:clock, Multiplier18:clock, Multiplier19:clock, Multiplier1:clock, Multiplier20:clock, Multiplier21:clock, Multiplier22:clock, Multiplier23:clock, Multiplier24:clock, Multiplier2:clock, Multiplier3:clock, Multiplier4:clock, Multiplier5:clock, Multiplier6:clock, Multiplier7:clock, Multiplier8:clock, Multiplier9:clock, Multiplier:clock, Parallel_Adder_Subtractor:clock, Pipelined_Adder:clock, Round:clk]
	signal clock_0_clock_output_reset                        : std_logic;                     -- Clock_0:aclr_out -> [Bus_Concatenation1:aclr, Bus_Concatenation:aclr, Memory_Delay:aclr, Multiplier10:aclr, Multiplier11:aclr, Multiplier12:aclr, Multiplier13:aclr, Multiplier14:aclr, Multiplier15:aclr, Multiplier16:aclr, Multiplier17:aclr, Multiplier18:aclr, Multiplier19:aclr, Multiplier1:aclr, Multiplier20:aclr, Multiplier21:aclr, Multiplier22:aclr, Multiplier23:aclr, Multiplier24:aclr, Multiplier2:aclr, Multiplier3:aclr, Multiplier4:aclr, Multiplier5:aclr, Multiplier6:aclr, Multiplier7:aclr, Multiplier8:aclr, Multiplier9:aclr, Multiplier:aclr, Parallel_Adder_Subtractor:aclr, Pipelined_Adder:aclr, Round:reset]

begin

	clock_0 : component alt_dspbuilder_clock_GNQFU4PUDH
		port map (
			clock_out => clock_0_clock_output_clk,   -- clock_output.clk
			aclr_out  => clock_0_clock_output_reset, --             .reset
			clock     => Clock,                      --        clock.clk
			aclr      => reset                       --             .reset
		);

	multiplier2 : component alt_dspbuilder_multiplier_GNNIEJHQ5V
		generic map (
			aWidth                         => 8,
			Signed                         => 0,
			bWidth                         => 26,
			DEDICATED_MULTIPLIER_CIRCUITRY => "NO",
			pipeline                       => 8,
			OutputLsb                      => 0,
			OutputMsb                      => 25
		)
		port map (
			clock     => clock_0_clock_output_clk,            -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,          --           .reset
			dataa     => data_02_0_output_wire,               --      dataa.wire
			datab     => constant2_output_wire,               --      datab.wire
			result    => multiplier2_result_wire,             --     result.wire
			user_aclr => multiplier2user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => clken_0_output_wire                  --        ena.wire
		);

	multiplier2user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplier2user_aclrgnd_output_wire  -- output.wire
		);

	multiplier1 : component alt_dspbuilder_multiplier_GNNIEJHQ5V
		generic map (
			aWidth                         => 8,
			Signed                         => 0,
			bWidth                         => 26,
			DEDICATED_MULTIPLIER_CIRCUITRY => "NO",
			pipeline                       => 8,
			OutputLsb                      => 0,
			OutputMsb                      => 25
		)
		port map (
			clock     => clock_0_clock_output_clk,            -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,          --           .reset
			dataa     => data_01_0_output_wire,               --      dataa.wire
			datab     => constant1_output_wire,               --      datab.wire
			result    => multiplier1_result_wire,             --     result.wire
			user_aclr => multiplier1user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => clken_0_output_wire                  --        ena.wire
		);

	multiplier1user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplier1user_aclrgnd_output_wire  -- output.wire
		);

	multiplier18 : component alt_dspbuilder_multiplier_GNNIEJHQ5V
		generic map (
			aWidth                         => 8,
			Signed                         => 0,
			bWidth                         => 26,
			DEDICATED_MULTIPLIER_CIRCUITRY => "NO",
			pipeline                       => 8,
			OutputLsb                      => 0,
			OutputMsb                      => 25
		)
		port map (
			clock     => clock_0_clock_output_clk,             -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,           --           .reset
			dataa     => data_33_0_output_wire,                --      dataa.wire
			datab     => constant18_output_wire,               --      datab.wire
			result    => multiplier18_result_wire,             --     result.wire
			user_aclr => multiplier18user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => clken_0_output_wire                   --        ena.wire
		);

	multiplier18user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplier18user_aclrgnd_output_wire  -- output.wire
		);

	multiplier4 : component alt_dspbuilder_multiplier_GNNIEJHQ5V
		generic map (
			aWidth                         => 8,
			Signed                         => 0,
			bWidth                         => 26,
			DEDICATED_MULTIPLIER_CIRCUITRY => "NO",
			pipeline                       => 8,
			OutputLsb                      => 0,
			OutputMsb                      => 25
		)
		port map (
			clock     => clock_0_clock_output_clk,            -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,          --           .reset
			dataa     => data_04_0_output_wire,               --      dataa.wire
			datab     => constant4_output_wire,               --      datab.wire
			result    => multiplier4_result_wire,             --     result.wire
			user_aclr => multiplier4user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => clken_0_output_wire                  --        ena.wire
		);

	multiplier4user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplier4user_aclrgnd_output_wire  -- output.wire
		);

	multiplier19 : component alt_dspbuilder_multiplier_GNNIEJHQ5V
		generic map (
			aWidth                         => 8,
			Signed                         => 0,
			bWidth                         => 26,
			DEDICATED_MULTIPLIER_CIRCUITRY => "NO",
			pipeline                       => 8,
			OutputLsb                      => 0,
			OutputMsb                      => 25
		)
		port map (
			clock     => clock_0_clock_output_clk,             -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,           --           .reset
			dataa     => data_34_0_output_wire,                --      dataa.wire
			datab     => constant19_output_wire,               --      datab.wire
			result    => multiplier19_result_wire,             --     result.wire
			user_aclr => multiplier19user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => clken_0_output_wire                   --        ena.wire
		);

	multiplier19user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplier19user_aclrgnd_output_wire  -- output.wire
		);

	multiplier3 : component alt_dspbuilder_multiplier_GNNIEJHQ5V
		generic map (
			aWidth                         => 8,
			Signed                         => 0,
			bWidth                         => 26,
			DEDICATED_MULTIPLIER_CIRCUITRY => "NO",
			pipeline                       => 8,
			OutputLsb                      => 0,
			OutputMsb                      => 25
		)
		port map (
			clock     => clock_0_clock_output_clk,            -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,          --           .reset
			dataa     => data_03_0_output_wire,               --      dataa.wire
			datab     => constant3_output_wire,               --      datab.wire
			result    => multiplier3_result_wire,             --     result.wire
			user_aclr => multiplier3user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => clken_0_output_wire                  --        ena.wire
		);

	multiplier3user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplier3user_aclrgnd_output_wire  -- output.wire
		);

	multiplier6 : component alt_dspbuilder_multiplier_GNNIEJHQ5V
		generic map (
			aWidth                         => 8,
			Signed                         => 0,
			bWidth                         => 26,
			DEDICATED_MULTIPLIER_CIRCUITRY => "NO",
			pipeline                       => 8,
			OutputLsb                      => 0,
			OutputMsb                      => 25
		)
		port map (
			clock     => clock_0_clock_output_clk,            -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,          --           .reset
			dataa     => data_11_0_output_wire,               --      dataa.wire
			datab     => constant6_output_wire,               --      datab.wire
			result    => multiplier6_result_wire,             --     result.wire
			user_aclr => multiplier6user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => clken_0_output_wire                  --        ena.wire
		);

	multiplier6user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplier6user_aclrgnd_output_wire  -- output.wire
		);

	multiplier5 : component alt_dspbuilder_multiplier_GNNIEJHQ5V
		generic map (
			aWidth                         => 8,
			Signed                         => 0,
			bWidth                         => 26,
			DEDICATED_MULTIPLIER_CIRCUITRY => "NO",
			pipeline                       => 8,
			OutputLsb                      => 0,
			OutputMsb                      => 25
		)
		port map (
			clock     => clock_0_clock_output_clk,            -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,          --           .reset
			dataa     => data_10_0_output_wire,               --      dataa.wire
			datab     => constant5_output_wire,               --      datab.wire
			result    => multiplier5_result_wire,             --     result.wire
			user_aclr => multiplier5user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => clken_0_output_wire                  --        ena.wire
		);

	multiplier5user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplier5user_aclrgnd_output_wire  -- output.wire
		);

	multiplier8 : component alt_dspbuilder_multiplier_GNNIEJHQ5V
		generic map (
			aWidth                         => 8,
			Signed                         => 0,
			bWidth                         => 26,
			DEDICATED_MULTIPLIER_CIRCUITRY => "NO",
			pipeline                       => 8,
			OutputLsb                      => 0,
			OutputMsb                      => 25
		)
		port map (
			clock     => clock_0_clock_output_clk,            -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,          --           .reset
			dataa     => data_13_0_output_wire,               --      dataa.wire
			datab     => constant8_output_wire,               --      datab.wire
			result    => multiplier8_result_wire,             --     result.wire
			user_aclr => multiplier8user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => clken_0_output_wire                  --        ena.wire
		);

	multiplier8user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplier8user_aclrgnd_output_wire  -- output.wire
		);

	constant26 : component alt_dspbuilder_constant_GN6SFEINY6
		generic map (
			BitPattern => "00",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 2
		)
		port map (
			output => constant26_output_wire  -- output.wire
		);

	multiplier7 : component alt_dspbuilder_multiplier_GNNIEJHQ5V
		generic map (
			aWidth                         => 8,
			Signed                         => 0,
			bWidth                         => 26,
			DEDICATED_MULTIPLIER_CIRCUITRY => "NO",
			pipeline                       => 8,
			OutputLsb                      => 0,
			OutputMsb                      => 25
		)
		port map (
			clock     => clock_0_clock_output_clk,            -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,          --           .reset
			dataa     => data_12_0_output_wire,               --      dataa.wire
			datab     => constant7_output_wire,               --      datab.wire
			result    => multiplier7_result_wire,             --     result.wire
			user_aclr => multiplier7user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => clken_0_output_wire                  --        ena.wire
		);

	multiplier7user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplier7user_aclrgnd_output_wire  -- output.wire
		);

	constant25 : component alt_dspbuilder_constant_GN6SFEINY6
		generic map (
			BitPattern => "00",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 2
		)
		port map (
			output => constant25_output_wire  -- output.wire
		);

	multiplier12 : component alt_dspbuilder_multiplier_GNNIEJHQ5V
		generic map (
			aWidth                         => 8,
			Signed                         => 0,
			bWidth                         => 26,
			DEDICATED_MULTIPLIER_CIRCUITRY => "NO",
			pipeline                       => 8,
			OutputLsb                      => 0,
			OutputMsb                      => 25
		)
		port map (
			clock     => clock_0_clock_output_clk,             -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,           --           .reset
			dataa     => data_22_0_output_wire,                --      dataa.wire
			datab     => constant12_output_wire,               --      datab.wire
			result    => multiplier12_result_wire,             --     result.wire
			user_aclr => multiplier12user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => clken_0_output_wire                   --        ena.wire
		);

	multiplier12user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplier12user_aclrgnd_output_wire  -- output.wire
		);

	constant24 : component alt_dspbuilder_constant_GN2DUUMQHA
		generic map (
			BitPattern => "00000000000000010000000000",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 26
		)
		port map (
			output => constant24_output_wire  -- output.wire
		);

	multiplier13 : component alt_dspbuilder_multiplier_GNNIEJHQ5V
		generic map (
			aWidth                         => 8,
			Signed                         => 0,
			bWidth                         => 26,
			DEDICATED_MULTIPLIER_CIRCUITRY => "NO",
			pipeline                       => 8,
			OutputLsb                      => 0,
			OutputMsb                      => 25
		)
		port map (
			clock     => clock_0_clock_output_clk,             -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,           --           .reset
			dataa     => data_23_0_output_wire,                --      dataa.wire
			datab     => constant13_output_wire,               --      datab.wire
			result    => multiplier13_result_wire,             --     result.wire
			user_aclr => multiplier13user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => clken_0_output_wire                   --        ena.wire
		);

	multiplier13user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplier13user_aclrgnd_output_wire  -- output.wire
		);

	multiplier9 : component alt_dspbuilder_multiplier_GNNIEJHQ5V
		generic map (
			aWidth                         => 8,
			Signed                         => 0,
			bWidth                         => 26,
			DEDICATED_MULTIPLIER_CIRCUITRY => "NO",
			pipeline                       => 8,
			OutputLsb                      => 0,
			OutputMsb                      => 25
		)
		port map (
			clock     => clock_0_clock_output_clk,            -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,          --           .reset
			dataa     => data_14_0_output_wire,               --      dataa.wire
			datab     => constant9_output_wire,               --      datab.wire
			result    => multiplier9_result_wire,             --     result.wire
			user_aclr => multiplier9user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => clken_0_output_wire                  --        ena.wire
		);

	multiplier9user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplier9user_aclrgnd_output_wire  -- output.wire
		);

	constant23 : component alt_dspbuilder_constant_GN52UV6F2X
		generic map (
			BitPattern => "00000000000001000000000000",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 26
		)
		port map (
			output => constant23_output_wire  -- output.wire
		);

	multiplier10 : component alt_dspbuilder_multiplier_GNNIEJHQ5V
		generic map (
			aWidth                         => 8,
			Signed                         => 0,
			bWidth                         => 26,
			DEDICATED_MULTIPLIER_CIRCUITRY => "NO",
			pipeline                       => 8,
			OutputLsb                      => 0,
			OutputMsb                      => 25
		)
		port map (
			clock     => clock_0_clock_output_clk,             -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,           --           .reset
			dataa     => data_20_0_output_wire,                --      dataa.wire
			datab     => constant10_output_wire,               --      datab.wire
			result    => multiplier10_result_wire,             --     result.wire
			user_aclr => multiplier10user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => clken_0_output_wire                   --        ena.wire
		);

	multiplier10user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplier10user_aclrgnd_output_wire  -- output.wire
		);

	constant22 : component alt_dspbuilder_constant_GNBQQQV5ZM
		generic map (
			BitPattern => "00000000000001100000000000",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 26
		)
		port map (
			output => constant22_output_wire  -- output.wire
		);

	multiplier11 : component alt_dspbuilder_multiplier_GNNIEJHQ5V
		generic map (
			aWidth                         => 8,
			Signed                         => 0,
			bWidth                         => 26,
			DEDICATED_MULTIPLIER_CIRCUITRY => "NO",
			pipeline                       => 8,
			OutputLsb                      => 0,
			OutputMsb                      => 25
		)
		port map (
			clock     => clock_0_clock_output_clk,             -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,           --           .reset
			dataa     => data_21_0_output_wire,                --      dataa.wire
			datab     => constant11_output_wire,               --      datab.wire
			result    => multiplier11_result_wire,             --     result.wire
			user_aclr => multiplier11user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => clken_0_output_wire                   --        ena.wire
		);

	multiplier11user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplier11user_aclrgnd_output_wire  -- output.wire
		);

	constant21 : component alt_dspbuilder_constant_GN52UV6F2X
		generic map (
			BitPattern => "00000000000001000000000000",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 26
		)
		port map (
			output => constant21_output_wire  -- output.wire
		);

	multiplier16 : component alt_dspbuilder_multiplier_GNNIEJHQ5V
		generic map (
			aWidth                         => 8,
			Signed                         => 0,
			bWidth                         => 26,
			DEDICATED_MULTIPLIER_CIRCUITRY => "NO",
			pipeline                       => 8,
			OutputLsb                      => 0,
			OutputMsb                      => 25
		)
		port map (
			clock     => clock_0_clock_output_clk,             -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,           --           .reset
			dataa     => data_31_0_output_wire,                --      dataa.wire
			datab     => constant16_output_wire,               --      datab.wire
			result    => multiplier16_result_wire,             --     result.wire
			user_aclr => multiplier16user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => clken_0_output_wire                   --        ena.wire
		);

	multiplier16user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplier16user_aclrgnd_output_wire  -- output.wire
		);

	constant20 : component alt_dspbuilder_constant_GN2DUUMQHA
		generic map (
			BitPattern => "00000000000000010000000000",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 26
		)
		port map (
			output => constant20_output_wire  -- output.wire
		);

	multiplier17 : component alt_dspbuilder_multiplier_GNNIEJHQ5V
		generic map (
			aWidth                         => 8,
			Signed                         => 0,
			bWidth                         => 26,
			DEDICATED_MULTIPLIER_CIRCUITRY => "NO",
			pipeline                       => 8,
			OutputLsb                      => 0,
			OutputMsb                      => 25
		)
		port map (
			clock     => clock_0_clock_output_clk,             -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,           --           .reset
			dataa     => data_32_0_output_wire,                --      dataa.wire
			datab     => constant17_output_wire,               --      datab.wire
			result    => multiplier17_result_wire,             --     result.wire
			user_aclr => multiplier17user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => clken_0_output_wire                   --        ena.wire
		);

	multiplier17user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplier17user_aclrgnd_output_wire  -- output.wire
		);

	multiplier14 : component alt_dspbuilder_multiplier_GNNIEJHQ5V
		generic map (
			aWidth                         => 8,
			Signed                         => 0,
			bWidth                         => 26,
			DEDICATED_MULTIPLIER_CIRCUITRY => "NO",
			pipeline                       => 8,
			OutputLsb                      => 0,
			OutputMsb                      => 25
		)
		port map (
			clock     => clock_0_clock_output_clk,             -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,           --           .reset
			dataa     => data_24_0_output_wire,                --      dataa.wire
			datab     => constant14_output_wire,               --      datab.wire
			result    => multiplier14_result_wire,             --     result.wire
			user_aclr => multiplier14user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => clken_0_output_wire                   --        ena.wire
		);

	multiplier14user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplier14user_aclrgnd_output_wire  -- output.wire
		);

	multiplier15 : component alt_dspbuilder_multiplier_GNNIEJHQ5V
		generic map (
			aWidth                         => 8,
			Signed                         => 0,
			bWidth                         => 26,
			DEDICATED_MULTIPLIER_CIRCUITRY => "NO",
			pipeline                       => 8,
			OutputLsb                      => 0,
			OutputMsb                      => 25
		)
		port map (
			clock     => clock_0_clock_output_clk,             -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,           --           .reset
			dataa     => data_30_0_output_wire,                --      dataa.wire
			datab     => constant15_output_wire,               --      datab.wire
			result    => multiplier15_result_wire,             --     result.wire
			user_aclr => multiplier15user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => clken_0_output_wire                   --        ena.wire
		);

	multiplier15user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplier15user_aclrgnd_output_wire  -- output.wire
		);

	data_33_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => data_33,               --  input.wire
			output => data_33_0_output_wire  -- output.wire
		);

	data_32_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => data_32,               --  input.wire
			output => data_32_0_output_wire  -- output.wire
		);

	data_34_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => data_34,               --  input.wire
			output => data_34_0_output_wire  -- output.wire
		);

	multiplier20 : component alt_dspbuilder_multiplier_GNNIEJHQ5V
		generic map (
			aWidth                         => 8,
			Signed                         => 0,
			bWidth                         => 26,
			DEDICATED_MULTIPLIER_CIRCUITRY => "NO",
			pipeline                       => 8,
			OutputLsb                      => 0,
			OutputMsb                      => 25
		)
		port map (
			clock     => clock_0_clock_output_clk,             -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,           --           .reset
			dataa     => data_40_0_output_wire,                --      dataa.wire
			datab     => constant20_output_wire,               --      datab.wire
			result    => multiplier20_result_wire,             --     result.wire
			user_aclr => multiplier20user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => clken_0_output_wire                   --        ena.wire
		);

	multiplier20user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplier20user_aclrgnd_output_wire  -- output.wire
		);

	data_31_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => data_31,               --  input.wire
			output => data_31_0_output_wire  -- output.wire
		);

	data_30_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => data_30,               --  input.wire
			output => data_30_0_output_wire  -- output.wire
		);

	constant2 : component alt_dspbuilder_constant_GNBQQQV5ZM
		generic map (
			BitPattern => "00000000000001100000000000",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 26
		)
		port map (
			output => constant2_output_wire  -- output.wire
		);

	multiplier23 : component alt_dspbuilder_multiplier_GNNIEJHQ5V
		generic map (
			aWidth                         => 8,
			Signed                         => 0,
			bWidth                         => 26,
			DEDICATED_MULTIPLIER_CIRCUITRY => "NO",
			pipeline                       => 8,
			OutputLsb                      => 0,
			OutputMsb                      => 25
		)
		port map (
			clock     => clock_0_clock_output_clk,             -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,           --           .reset
			dataa     => data_43_0_output_wire,                --      dataa.wire
			datab     => constant23_output_wire,               --      datab.wire
			result    => multiplier23_result_wire,             --     result.wire
			user_aclr => multiplier23user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => clken_0_output_wire                   --        ena.wire
		);

	multiplier23user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplier23user_aclrgnd_output_wire  -- output.wire
		);

	constant3 : component alt_dspbuilder_constant_GN52UV6F2X
		generic map (
			BitPattern => "00000000000001000000000000",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 26
		)
		port map (
			output => constant3_output_wire  -- output.wire
		);

	multiplier24 : component alt_dspbuilder_multiplier_GNNIEJHQ5V
		generic map (
			aWidth                         => 8,
			Signed                         => 0,
			bWidth                         => 26,
			DEDICATED_MULTIPLIER_CIRCUITRY => "NO",
			pipeline                       => 8,
			OutputLsb                      => 0,
			OutputMsb                      => 25
		)
		port map (
			clock     => clock_0_clock_output_clk,             -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,           --           .reset
			dataa     => data_44_0_output_wire,                --      dataa.wire
			datab     => constant24_output_wire,               --      datab.wire
			result    => multiplier24_result_wire,             --     result.wire
			user_aclr => multiplier24user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => clken_0_output_wire                   --        ena.wire
		);

	multiplier24user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplier24user_aclrgnd_output_wire  -- output.wire
		);

	multiplier21 : component alt_dspbuilder_multiplier_GNNIEJHQ5V
		generic map (
			aWidth                         => 8,
			Signed                         => 0,
			bWidth                         => 26,
			DEDICATED_MULTIPLIER_CIRCUITRY => "NO",
			pipeline                       => 8,
			OutputLsb                      => 0,
			OutputMsb                      => 25
		)
		port map (
			clock     => clock_0_clock_output_clk,             -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,           --           .reset
			dataa     => data_41_0_output_wire,                --      dataa.wire
			datab     => constant21_output_wire,               --      datab.wire
			result    => multiplier21_result_wire,             --     result.wire
			user_aclr => multiplier21user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => clken_0_output_wire                   --        ena.wire
		);

	multiplier21user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplier21user_aclrgnd_output_wire  -- output.wire
		);

	constant1 : component alt_dspbuilder_constant_GN52UV6F2X
		generic map (
			BitPattern => "00000000000001000000000000",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 26
		)
		port map (
			output => constant1_output_wire  -- output.wire
		);

	multiplier22 : component alt_dspbuilder_multiplier_GNNIEJHQ5V
		generic map (
			aWidth                         => 8,
			Signed                         => 0,
			bWidth                         => 26,
			DEDICATED_MULTIPLIER_CIRCUITRY => "NO",
			pipeline                       => 8,
			OutputLsb                      => 0,
			OutputMsb                      => 25
		)
		port map (
			clock     => clock_0_clock_output_clk,             -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,           --           .reset
			dataa     => data_42_0_output_wire,                --      dataa.wire
			datab     => constant22_output_wire,               --      datab.wire
			result    => multiplier22_result_wire,             --     result.wire
			user_aclr => multiplier22user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => clken_0_output_wire                   --        ena.wire
		);

	multiplier22user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplier22user_aclrgnd_output_wire  -- output.wire
		);

	data_00_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => data_00,               --  input.wire
			output => data_00_0_output_wire  -- output.wire
		);

	data_44_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => data_44,               --  input.wire
			output => data_44_0_output_wire  -- output.wire
		);

	bus_concatenation1 : component alt_dspbuilder_bus_concat_GNKLOJ6ING
		generic map (
			widthA => 2,
			widthB => 8
		)
		port map (
			clock  => clock_0_clock_output_clk,       -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,     --           .reset
			a      => constant25_output_wire,         --          a.wire
			b      => cast0_output_wire,              --          b.wire
			output => bus_concatenation1_output_wire  --     output.wire
		);

	data_43_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => data_43,               --  input.wire
			output => data_43_0_output_wire  -- output.wire
		);

	data_02_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => data_02,               --  input.wire
			output => data_02_0_output_wire  -- output.wire
		);

	constant8 : component alt_dspbuilder_constant_GN42V6LR6J
		generic map (
			BitPattern => "00000000000100000000000000",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 26
		)
		port map (
			output => constant8_output_wire  -- output.wire
		);

	data_01_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => data_01,               --  input.wire
			output => data_01_0_output_wire  -- output.wire
		);

	constant9 : component alt_dspbuilder_constant_GN52UV6F2X
		generic map (
			BitPattern => "00000000000001000000000000",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 26
		)
		port map (
			output => constant9_output_wire  -- output.wire
		);

	data_40_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => data_40,               --  input.wire
			output => data_40_0_output_wire  -- output.wire
		);

	constant6 : component alt_dspbuilder_constant_GN42V6LR6J
		generic map (
			BitPattern => "00000000000100000000000000",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 26
		)
		port map (
			output => constant6_output_wire  -- output.wire
		);

	constant7 : component alt_dspbuilder_constant_GN3UR3AYSK
		generic map (
			BitPattern => "00000000000110000000000000",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 26
		)
		port map (
			output => constant7_output_wire  -- output.wire
		);

	data_42_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => data_42,               --  input.wire
			output => data_42_0_output_wire  -- output.wire
		);

	constant4 : component alt_dspbuilder_constant_GN2DUUMQHA
		generic map (
			BitPattern => "00000000000000010000000000",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 26
		)
		port map (
			output => constant4_output_wire  -- output.wire
		);

	data_41_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => data_41,               --  input.wire
			output => data_41_0_output_wire  -- output.wire
		);

	constant5 : component alt_dspbuilder_constant_GN52UV6F2X
		generic map (
			BitPattern => "00000000000001000000000000",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 26
		)
		port map (
			output => constant5_output_wire  -- output.wire
		);

	pixel_out_0 : component alt_dspbuilder_port_GNEPKLLZKY
		port map (
			input  => parallel_adder_subtractor_result_wire, --  input.wire
			output => pixel_out                              -- output.wire
		);

	data_04_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => data_04,               --  input.wire
			output => data_04_0_output_wire  -- output.wire
		);

	data_03_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => data_03,               --  input.wire
			output => data_03_0_output_wire  -- output.wire
		);

	bus_concatenation : component alt_dspbuilder_bus_concat_GNKLOJ6ING
		generic map (
			widthA => 2,
			widthB => 8
		)
		port map (
			clock  => clock_0_clock_output_clk,      -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,    --           .reset
			a      => constant26_output_wire,        --          a.wire
			b      => cast27_output_wire,            --          b.wire
			output => bus_concatenation_output_wire  --     output.wire
		);

	pipelined_adder : component alt_dspbuilder_pipelined_adder_GNY2JEH574
		generic map (
			pipeline => 1,
			width    => 10
		)
		port map (
			clock     => clock_0_clock_output_clk,                -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,              --           .reset
			dataa     => bus_concatenation1_output_wire,          --      dataa.wire
			datab     => bus_concatenation_output_wire,           --      datab.wire
			result    => pipelined_adder_result_wire,             --     result.wire
			user_aclr => pipelined_adderuser_aclrgnd_output_wire, --  user_aclr.wire
			ena       => clken_0_output_wire                      --        ena.wire
		);

	pipelined_adderuser_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => pipelined_adderuser_aclrgnd_output_wire  -- output.wire
		);

	data_11_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => data_11,               --  input.wire
			output => data_11_0_output_wire  -- output.wire
		);

	data_10_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => data_10,               --  input.wire
			output => data_10_0_output_wire  -- output.wire
		);

	data_13_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => data_13,               --  input.wire
			output => data_13_0_output_wire  -- output.wire
		);

	data_12_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => data_12,               --  input.wire
			output => data_12_0_output_wire  -- output.wire
		);

	pixel_diff_0 : component alt_dspbuilder_port_GNSSYS4J5R
		port map (
			input  => pipelined_adder_result_wire, --  input.wire
			output => pixel_diff                   -- output.wire
		);

	multiplier : component alt_dspbuilder_multiplier_GNNIEJHQ5V
		generic map (
			aWidth                         => 8,
			Signed                         => 0,
			bWidth                         => 26,
			DEDICATED_MULTIPLIER_CIRCUITRY => "NO",
			pipeline                       => 8,
			OutputLsb                      => 0,
			OutputMsb                      => 25
		)
		port map (
			clock     => clock_0_clock_output_clk,           -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,         --           .reset
			dataa     => data_00_0_output_wire,              --      dataa.wire
			datab     => constant_1_output_wire,             --      datab.wire
			result    => multiplier_result_wire,             --     result.wire
			user_aclr => multiplieruser_aclrgnd_output_wire, --  user_aclr.wire
			ena       => clken_0_output_wire                 --        ena.wire
		);

	multiplieruser_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplieruser_aclrgnd_output_wire  -- output.wire
		);

	round : component alt_dspbuilder_round_GNWBUVGWWO
		generic map (
			OUT_WIDTH_g     => 8,
			IN_WIDTH_g      => 26,
			PIPELINE_g      => 0,
			ROUNDING_TYPE_g => "ROUND_UP",
			SIGNED_g        => 0
		)
		port map (
			clk       => clock_0_clock_output_clk,      -- clk_reset.clk
			reset     => clock_0_clock_output_reset,    --          .reset
			datain    => cast26_output_wire,            --    datain.wire
			dataout   => round_dataout_wire,            --   dataout.wire
			ena       => roundenavcc_output_wire,       --       ena.wire
			user_aclr => rounduser_aclrgnd_output_wire  -- user_aclr.wire
		);

	rounduser_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => rounduser_aclrgnd_output_wire  -- output.wire
		);

	roundenavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => roundenavcc_output_wire  -- output.wire
		);

	roundresetgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => roundresetgnd_output_wire  -- output.wire
		);

	data_14_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => data_14,               --  input.wire
			output => data_14_0_output_wire  -- output.wire
		);

	constant19 : component alt_dspbuilder_constant_GN52UV6F2X
		generic map (
			BitPattern => "00000000000001000000000000",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 26
		)
		port map (
			output => constant19_output_wire  -- output.wire
		);

	constant18 : component alt_dspbuilder_constant_GN42V6LR6J
		generic map (
			BitPattern => "00000000000100000000000000",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 26
		)
		port map (
			output => constant18_output_wire  -- output.wire
		);

	parallel_adder_subtractor : component alt_dspbuilder_parallel_adder_GN5CSCONM5
		generic map (
			dataWidth     => 27,
			direction     => "+",
			MaskValue     => "1",
			pipeline      => 1,
			number_inputs => 25
		)
		port map (
			clock     => clock_0_clock_output_clk,                          -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,                        --           .reset
			result    => parallel_adder_subtractor_result_wire,             --     result.wire
			user_aclr => parallel_adder_subtractoruser_aclrgnd_output_wire, --  user_aclr.wire
			ena       => clken_0_output_wire,                               --        ena.wire
			data0     => cast1_output_wire,                                 --      data0.wire
			data1     => cast2_output_wire,                                 --      data1.wire
			data2     => cast3_output_wire,                                 --      data2.wire
			data3     => cast4_output_wire,                                 --      data3.wire
			data4     => cast5_output_wire,                                 --      data4.wire
			data5     => cast6_output_wire,                                 --      data5.wire
			data6     => cast7_output_wire,                                 --      data6.wire
			data7     => cast8_output_wire,                                 --      data7.wire
			data8     => cast9_output_wire,                                 --      data8.wire
			data9     => cast10_output_wire,                                --      data9.wire
			data10    => cast11_output_wire,                                --     data10.wire
			data11    => cast12_output_wire,                                --     data11.wire
			data12    => cast13_output_wire,                                --     data12.wire
			data13    => cast14_output_wire,                                --     data13.wire
			data14    => cast15_output_wire,                                --     data14.wire
			data15    => cast16_output_wire,                                --     data15.wire
			data16    => cast17_output_wire,                                --     data16.wire
			data17    => cast18_output_wire,                                --     data17.wire
			data18    => cast19_output_wire,                                --     data18.wire
			data19    => cast20_output_wire,                                --     data19.wire
			data20    => cast21_output_wire,                                --     data20.wire
			data21    => cast22_output_wire,                                --     data21.wire
			data22    => cast23_output_wire,                                --     data22.wire
			data23    => cast24_output_wire,                                --     data23.wire
			data24    => cast25_output_wire                                 --     data24.wire
		);

	parallel_adder_subtractoruser_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => parallel_adder_subtractoruser_aclrgnd_output_wire  -- output.wire
		);

	constant17 : component alt_dspbuilder_constant_GN3UR3AYSK
		generic map (
			BitPattern => "00000000000110000000000000",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 26
		)
		port map (
			output => constant17_output_wire  -- output.wire
		);

	constant16 : component alt_dspbuilder_constant_GN42V6LR6J
		generic map (
			BitPattern => "00000000000100000000000000",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 26
		)
		port map (
			output => constant16_output_wire  -- output.wire
		);

	constant15 : component alt_dspbuilder_constant_GN52UV6F2X
		generic map (
			BitPattern => "00000000000001000000000000",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 26
		)
		port map (
			output => constant15_output_wire  -- output.wire
		);

	constant14 : component alt_dspbuilder_constant_GNBQQQV5ZM
		generic map (
			BitPattern => "00000000000001100000000000",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 26
		)
		port map (
			output => constant14_output_wire  -- output.wire
		);

	constant13 : component alt_dspbuilder_constant_GN3UR3AYSK
		generic map (
			BitPattern => "00000000000110000000000000",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 26
		)
		port map (
			output => constant13_output_wire  -- output.wire
		);

	constant12 : component alt_dspbuilder_constant_GNHUGKQYBA
		generic map (
			BitPattern => "00000000001001000000000000",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 26
		)
		port map (
			output => constant12_output_wire  -- output.wire
		);

	constant11 : component alt_dspbuilder_constant_GN3UR3AYSK
		generic map (
			BitPattern => "00000000000110000000000000",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 26
		)
		port map (
			output => constant11_output_wire  -- output.wire
		);

	constant10 : component alt_dspbuilder_constant_GNBQQQV5ZM
		generic map (
			BitPattern => "00000000000001100000000000",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 26
		)
		port map (
			output => constant10_output_wire  -- output.wire
		);

	clken_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => clken,               --  input.wire
			output => clken_0_output_wire  -- output.wire
		);

	data_22_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => data_22,               --  input.wire
			output => data_22_0_output_wire  -- output.wire
		);

	data_21_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => data_21,               --  input.wire
			output => data_21_0_output_wire  -- output.wire
		);

	data_24_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => data_24,               --  input.wire
			output => data_24_0_output_wire  -- output.wire
		);

	data_23_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => data_23,               --  input.wire
			output => data_23_0_output_wire  -- output.wire
		);

	data_20_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => data_20,               --  input.wire
			output => data_20_0_output_wire  -- output.wire
		);

	constant_1 : component alt_dspbuilder_constant_GN2DUUMQHA
		generic map (
			BitPattern => "00000000000000010000000000",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 26
		)
		port map (
			output => constant_1_output_wire  -- output.wire
		);

	memory_delay : component alt_dspbuilder_memdelay_GND4ZY57YF
		generic map (
			RAMTYPE => "AUTO",
			WIDTH   => 8,
			DELAY   => 13
		)
		port map (
			clock     => clock_0_clock_output_clk,             -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,           --           .reset
			input     => data_22_0_output_wire,                --      input.wire
			output    => memory_delay_output_wire,             --     output.wire
			user_aclr => memory_delayuser_aclrgnd_output_wire, --  user_aclr.wire
			ena       => clken_0_output_wire                   --        ena.wire
		);

	memory_delayuser_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => memory_delayuser_aclrgnd_output_wire  -- output.wire
		);

	cast0 : component alt_dspbuilder_cast_GNBZR5PMEK
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => memory_delay_output_wire, --  input.wire
			output => cast0_output_wire         -- output.wire
		);

	cast1 : component alt_dspbuilder_cast_GNMLNX2RCD
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => multiplier_result_wire, --  input.wire
			output => cast1_output_wire       -- output.wire
		);

	cast2 : component alt_dspbuilder_cast_GNMLNX2RCD
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => multiplier1_result_wire, --  input.wire
			output => cast2_output_wire        -- output.wire
		);

	cast3 : component alt_dspbuilder_cast_GNMLNX2RCD
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => multiplier2_result_wire, --  input.wire
			output => cast3_output_wire        -- output.wire
		);

	cast4 : component alt_dspbuilder_cast_GNMLNX2RCD
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => multiplier3_result_wire, --  input.wire
			output => cast4_output_wire        -- output.wire
		);

	cast5 : component alt_dspbuilder_cast_GNMLNX2RCD
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => multiplier4_result_wire, --  input.wire
			output => cast5_output_wire        -- output.wire
		);

	cast6 : component alt_dspbuilder_cast_GNMLNX2RCD
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => multiplier5_result_wire, --  input.wire
			output => cast6_output_wire        -- output.wire
		);

	cast7 : component alt_dspbuilder_cast_GNMLNX2RCD
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => multiplier6_result_wire, --  input.wire
			output => cast7_output_wire        -- output.wire
		);

	cast8 : component alt_dspbuilder_cast_GNMLNX2RCD
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => multiplier7_result_wire, --  input.wire
			output => cast8_output_wire        -- output.wire
		);

	cast9 : component alt_dspbuilder_cast_GNMLNX2RCD
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => multiplier8_result_wire, --  input.wire
			output => cast9_output_wire        -- output.wire
		);

	cast10 : component alt_dspbuilder_cast_GNMLNX2RCD
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => multiplier9_result_wire, --  input.wire
			output => cast10_output_wire       -- output.wire
		);

	cast11 : component alt_dspbuilder_cast_GNMLNX2RCD
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => multiplier10_result_wire, --  input.wire
			output => cast11_output_wire        -- output.wire
		);

	cast12 : component alt_dspbuilder_cast_GNMLNX2RCD
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => multiplier11_result_wire, --  input.wire
			output => cast12_output_wire        -- output.wire
		);

	cast13 : component alt_dspbuilder_cast_GNMLNX2RCD
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => multiplier12_result_wire, --  input.wire
			output => cast13_output_wire        -- output.wire
		);

	cast14 : component alt_dspbuilder_cast_GNMLNX2RCD
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => multiplier13_result_wire, --  input.wire
			output => cast14_output_wire        -- output.wire
		);

	cast15 : component alt_dspbuilder_cast_GNMLNX2RCD
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => multiplier14_result_wire, --  input.wire
			output => cast15_output_wire        -- output.wire
		);

	cast16 : component alt_dspbuilder_cast_GNMLNX2RCD
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => multiplier15_result_wire, --  input.wire
			output => cast16_output_wire        -- output.wire
		);

	cast17 : component alt_dspbuilder_cast_GNMLNX2RCD
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => multiplier16_result_wire, --  input.wire
			output => cast17_output_wire        -- output.wire
		);

	cast18 : component alt_dspbuilder_cast_GNMLNX2RCD
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => multiplier17_result_wire, --  input.wire
			output => cast18_output_wire        -- output.wire
		);

	cast19 : component alt_dspbuilder_cast_GNMLNX2RCD
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => multiplier18_result_wire, --  input.wire
			output => cast19_output_wire        -- output.wire
		);

	cast20 : component alt_dspbuilder_cast_GNMLNX2RCD
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => multiplier19_result_wire, --  input.wire
			output => cast20_output_wire        -- output.wire
		);

	cast21 : component alt_dspbuilder_cast_GNMLNX2RCD
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => multiplier20_result_wire, --  input.wire
			output => cast21_output_wire        -- output.wire
		);

	cast22 : component alt_dspbuilder_cast_GNMLNX2RCD
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => multiplier21_result_wire, --  input.wire
			output => cast22_output_wire        -- output.wire
		);

	cast23 : component alt_dspbuilder_cast_GNMLNX2RCD
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => multiplier22_result_wire, --  input.wire
			output => cast23_output_wire        -- output.wire
		);

	cast24 : component alt_dspbuilder_cast_GNMLNX2RCD
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => multiplier23_result_wire, --  input.wire
			output => cast24_output_wire        -- output.wire
		);

	cast25 : component alt_dspbuilder_cast_GNMLNX2RCD
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => multiplier24_result_wire, --  input.wire
			output => cast25_output_wire        -- output.wire
		);

	cast26 : component alt_dspbuilder_cast_GNHYNEPC7U
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => parallel_adder_subtractor_result_wire, --  input.wire
			output => cast26_output_wire                     -- output.wire
		);

	cast27 : component alt_dspbuilder_cast_GNBZR5PMEK
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => round_dataout_wire, --  input.wire
			output => cast27_output_wire  -- output.wire
		);

end architecture rtl; -- of gaussian_ip_GN_gaussian_ip_Fusion_Decomposition_3_multiplier_accumulator
