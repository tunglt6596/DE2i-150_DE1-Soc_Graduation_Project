// Computer_System.v

// Generated using ACDS version 17.1 590

`timescale 1 ps / 1 ps
module Computer_System (
		output wire        hps_io_hps_io_emac1_inst_TX_CLK, //               hps_io.hps_io_emac1_inst_TX_CLK
		output wire        hps_io_hps_io_emac1_inst_TXD0,   //                     .hps_io_emac1_inst_TXD0
		output wire        hps_io_hps_io_emac1_inst_TXD1,   //                     .hps_io_emac1_inst_TXD1
		output wire        hps_io_hps_io_emac1_inst_TXD2,   //                     .hps_io_emac1_inst_TXD2
		output wire        hps_io_hps_io_emac1_inst_TXD3,   //                     .hps_io_emac1_inst_TXD3
		input  wire        hps_io_hps_io_emac1_inst_RXD0,   //                     .hps_io_emac1_inst_RXD0
		inout  wire        hps_io_hps_io_emac1_inst_MDIO,   //                     .hps_io_emac1_inst_MDIO
		output wire        hps_io_hps_io_emac1_inst_MDC,    //                     .hps_io_emac1_inst_MDC
		input  wire        hps_io_hps_io_emac1_inst_RX_CTL, //                     .hps_io_emac1_inst_RX_CTL
		output wire        hps_io_hps_io_emac1_inst_TX_CTL, //                     .hps_io_emac1_inst_TX_CTL
		input  wire        hps_io_hps_io_emac1_inst_RX_CLK, //                     .hps_io_emac1_inst_RX_CLK
		input  wire        hps_io_hps_io_emac1_inst_RXD1,   //                     .hps_io_emac1_inst_RXD1
		input  wire        hps_io_hps_io_emac1_inst_RXD2,   //                     .hps_io_emac1_inst_RXD2
		input  wire        hps_io_hps_io_emac1_inst_RXD3,   //                     .hps_io_emac1_inst_RXD3
		inout  wire        hps_io_hps_io_qspi_inst_IO0,     //                     .hps_io_qspi_inst_IO0
		inout  wire        hps_io_hps_io_qspi_inst_IO1,     //                     .hps_io_qspi_inst_IO1
		inout  wire        hps_io_hps_io_qspi_inst_IO2,     //                     .hps_io_qspi_inst_IO2
		inout  wire        hps_io_hps_io_qspi_inst_IO3,     //                     .hps_io_qspi_inst_IO3
		output wire        hps_io_hps_io_qspi_inst_SS0,     //                     .hps_io_qspi_inst_SS0
		output wire        hps_io_hps_io_qspi_inst_CLK,     //                     .hps_io_qspi_inst_CLK
		inout  wire        hps_io_hps_io_sdio_inst_CMD,     //                     .hps_io_sdio_inst_CMD
		inout  wire        hps_io_hps_io_sdio_inst_D0,      //                     .hps_io_sdio_inst_D0
		inout  wire        hps_io_hps_io_sdio_inst_D1,      //                     .hps_io_sdio_inst_D1
		output wire        hps_io_hps_io_sdio_inst_CLK,     //                     .hps_io_sdio_inst_CLK
		inout  wire        hps_io_hps_io_sdio_inst_D2,      //                     .hps_io_sdio_inst_D2
		inout  wire        hps_io_hps_io_sdio_inst_D3,      //                     .hps_io_sdio_inst_D3
		inout  wire        hps_io_hps_io_usb1_inst_D0,      //                     .hps_io_usb1_inst_D0
		inout  wire        hps_io_hps_io_usb1_inst_D1,      //                     .hps_io_usb1_inst_D1
		inout  wire        hps_io_hps_io_usb1_inst_D2,      //                     .hps_io_usb1_inst_D2
		inout  wire        hps_io_hps_io_usb1_inst_D3,      //                     .hps_io_usb1_inst_D3
		inout  wire        hps_io_hps_io_usb1_inst_D4,      //                     .hps_io_usb1_inst_D4
		inout  wire        hps_io_hps_io_usb1_inst_D5,      //                     .hps_io_usb1_inst_D5
		inout  wire        hps_io_hps_io_usb1_inst_D6,      //                     .hps_io_usb1_inst_D6
		inout  wire        hps_io_hps_io_usb1_inst_D7,      //                     .hps_io_usb1_inst_D7
		input  wire        hps_io_hps_io_usb1_inst_CLK,     //                     .hps_io_usb1_inst_CLK
		output wire        hps_io_hps_io_usb1_inst_STP,     //                     .hps_io_usb1_inst_STP
		input  wire        hps_io_hps_io_usb1_inst_DIR,     //                     .hps_io_usb1_inst_DIR
		input  wire        hps_io_hps_io_usb1_inst_NXT,     //                     .hps_io_usb1_inst_NXT
		output wire        hps_io_hps_io_spim1_inst_CLK,    //                     .hps_io_spim1_inst_CLK
		output wire        hps_io_hps_io_spim1_inst_MOSI,   //                     .hps_io_spim1_inst_MOSI
		input  wire        hps_io_hps_io_spim1_inst_MISO,   //                     .hps_io_spim1_inst_MISO
		output wire        hps_io_hps_io_spim1_inst_SS0,    //                     .hps_io_spim1_inst_SS0
		input  wire        hps_io_hps_io_uart0_inst_RX,     //                     .hps_io_uart0_inst_RX
		output wire        hps_io_hps_io_uart0_inst_TX,     //                     .hps_io_uart0_inst_TX
		inout  wire        hps_io_hps_io_i2c0_inst_SDA,     //                     .hps_io_i2c0_inst_SDA
		inout  wire        hps_io_hps_io_i2c0_inst_SCL,     //                     .hps_io_i2c0_inst_SCL
		inout  wire        hps_io_hps_io_i2c1_inst_SDA,     //                     .hps_io_i2c1_inst_SDA
		inout  wire        hps_io_hps_io_i2c1_inst_SCL,     //                     .hps_io_i2c1_inst_SCL
		inout  wire        hps_io_hps_io_gpio_inst_GPIO09,  //                     .hps_io_gpio_inst_GPIO09
		inout  wire        hps_io_hps_io_gpio_inst_GPIO35,  //                     .hps_io_gpio_inst_GPIO35
		inout  wire        hps_io_hps_io_gpio_inst_GPIO40,  //                     .hps_io_gpio_inst_GPIO40
		inout  wire        hps_io_hps_io_gpio_inst_GPIO41,  //                     .hps_io_gpio_inst_GPIO41
		inout  wire        hps_io_hps_io_gpio_inst_GPIO48,  //                     .hps_io_gpio_inst_GPIO48
		inout  wire        hps_io_hps_io_gpio_inst_GPIO53,  //                     .hps_io_gpio_inst_GPIO53
		inout  wire        hps_io_hps_io_gpio_inst_GPIO54,  //                     .hps_io_gpio_inst_GPIO54
		inout  wire        hps_io_hps_io_gpio_inst_GPIO61,  //                     .hps_io_gpio_inst_GPIO61
		output wire [14:0] memory_mem_a,                    //               memory.mem_a
		output wire [2:0]  memory_mem_ba,                   //                     .mem_ba
		output wire        memory_mem_ck,                   //                     .mem_ck
		output wire        memory_mem_ck_n,                 //                     .mem_ck_n
		output wire        memory_mem_cke,                  //                     .mem_cke
		output wire        memory_mem_cs_n,                 //                     .mem_cs_n
		output wire        memory_mem_ras_n,                //                     .mem_ras_n
		output wire        memory_mem_cas_n,                //                     .mem_cas_n
		output wire        memory_mem_we_n,                 //                     .mem_we_n
		output wire        memory_mem_reset_n,              //                     .mem_reset_n
		inout  wire [31:0] memory_mem_dq,                   //                     .mem_dq
		inout  wire [3:0]  memory_mem_dqs,                  //                     .mem_dqs
		inout  wire [3:0]  memory_mem_dqs_n,                //                     .mem_dqs_n
		output wire        memory_mem_odt,                  //                     .mem_odt
		output wire [3:0]  memory_mem_dm,                   //                     .mem_dm
		input  wire        memory_oct_rzqin,                //                     .oct_rzqin
		input  wire        system_pll_ref_clk_clk,          //   system_pll_ref_clk.clk
		input  wire        system_pll_ref_reset_reset,      // system_pll_ref_reset.reset
		output wire        vga_CLK,                         //                  vga.CLK
		output wire        vga_HS,                          //                     .HS
		output wire        vga_VS,                          //                     .VS
		output wire        vga_BLANK,                       //                     .BLANK
		output wire        vga_SYNC,                        //                     .SYNC
		output wire [7:0]  vga_R,                           //                     .R
		output wire [7:0]  vga_G,                           //                     .G
		output wire [7:0]  vga_B,                           //                     .B
		output wire        vga_clk_clk,                     //              vga_clk.clk
		input  wire        vga_pll_ref_clk_clk,             //      vga_pll_ref_clk.clk
		input  wire        vga_pll_ref_reset_reset          //    vga_pll_ref_reset.reset
	);

	wire         padding_1_avalon_clipper_source_valid;                              // PADDING_1:stream_out_valid -> FUSION:sink1_valid
	wire   [7:0] padding_1_avalon_clipper_source_data;                               // PADDING_1:stream_out_data -> FUSION:sink1_data
	wire         padding_1_avalon_clipper_source_ready;                              // FUSION:sink1_ready -> PADDING_1:stream_out_ready
	wire         padding_1_avalon_clipper_source_startofpacket;                      // PADDING_1:stream_out_startofpacket -> FUSION:sink1_sop
	wire         padding_1_avalon_clipper_source_endofpacket;                        // PADDING_1:stream_out_endofpacket -> FUSION:sink1_eop
	wire         padding_2_avalon_clipper_source_valid;                              // PADDING_2:stream_out_valid -> FUSION:sink2_valid
	wire   [7:0] padding_2_avalon_clipper_source_data;                               // PADDING_2:stream_out_data -> FUSION:sink2_data
	wire         padding_2_avalon_clipper_source_ready;                              // FUSION:sink2_ready -> PADDING_2:stream_out_ready
	wire         padding_2_avalon_clipper_source_startofpacket;                      // PADDING_2:stream_out_startofpacket -> FUSION:sink2_sop
	wire         padding_2_avalon_clipper_source_endofpacket;                        // PADDING_2:stream_out_endofpacket -> FUSION:sink2_eop
	wire         dma_1_avalon_pixel_source_valid;                                    // DMA_1:stream_valid -> BUFFER_1:in_valid
	wire   [7:0] dma_1_avalon_pixel_source_data;                                     // DMA_1:stream_data -> BUFFER_1:in_data
	wire         dma_1_avalon_pixel_source_ready;                                    // BUFFER_1:in_ready -> DMA_1:stream_ready
	wire         dma_1_avalon_pixel_source_startofpacket;                            // DMA_1:stream_startofpacket -> BUFFER_1:in_startofpacket
	wire         dma_1_avalon_pixel_source_endofpacket;                              // DMA_1:stream_endofpacket -> BUFFER_1:in_endofpacket
	wire         dma_2_avalon_pixel_source_valid;                                    // DMA_2:stream_valid -> BUFFER_2:in_valid
	wire   [7:0] dma_2_avalon_pixel_source_data;                                     // DMA_2:stream_data -> BUFFER_2:in_data
	wire         dma_2_avalon_pixel_source_ready;                                    // BUFFER_2:in_ready -> DMA_2:stream_ready
	wire         dma_2_avalon_pixel_source_startofpacket;                            // DMA_2:stream_startofpacket -> BUFFER_2:in_startofpacket
	wire         dma_2_avalon_pixel_source_endofpacket;                              // DMA_2:stream_endofpacket -> BUFFER_2:in_endofpacket
	wire         fusion_data_source_valid;                                           // FUSION:source_valid -> DMA_WRITE:stream_valid
	wire   [7:0] fusion_data_source_data;                                            // FUSION:source_data -> DMA_WRITE:stream_data
	wire         fusion_data_source_ready;                                           // DMA_WRITE:stream_ready -> FUSION:source_ready
	wire         fusion_data_source_startofpacket;                                   // FUSION:source_sop -> DMA_WRITE:stream_startofpacket
	wire         fusion_data_source_endofpacket;                                     // FUSION:source_eop -> DMA_WRITE:stream_endofpacket
	wire         buffer_1_out_valid;                                                 // BUFFER_1:out_valid -> PADDING_1:stream_in_valid
	wire   [7:0] buffer_1_out_data;                                                  // BUFFER_1:out_data -> PADDING_1:stream_in_data
	wire         buffer_1_out_ready;                                                 // PADDING_1:stream_in_ready -> BUFFER_1:out_ready
	wire         buffer_1_out_startofpacket;                                         // BUFFER_1:out_startofpacket -> PADDING_1:stream_in_startofpacket
	wire         buffer_1_out_endofpacket;                                           // BUFFER_1:out_endofpacket -> PADDING_1:stream_in_endofpacket
	wire         buffer_2_out_valid;                                                 // BUFFER_2:out_valid -> PADDING_2:stream_in_valid
	wire   [7:0] buffer_2_out_data;                                                  // BUFFER_2:out_data -> PADDING_2:stream_in_data
	wire         buffer_2_out_ready;                                                 // PADDING_2:stream_in_ready -> BUFFER_2:out_ready
	wire         buffer_2_out_startofpacket;                                         // BUFFER_2:out_startofpacket -> PADDING_2:stream_in_startofpacket
	wire         buffer_2_out_endofpacket;                                           // BUFFER_2:out_endofpacket -> PADDING_2:stream_in_endofpacket
	wire         system_pll_sys_clk_clk;                                             // SYSTEM_PLL:sys_clk_clk -> [ARM_A9_HPS:f2h_axi_clk, ARM_A9_HPS:h2f_axi_clk, ARM_A9_HPS:h2f_lw_axi_clk, BUFFER_1:clk, BUFFER_2:clk, DMA_1:clk, DMA_2:clk, DMA_WRITE:clk, FUSION:Clock, PADDING_1:clk, PADDING_2:clk, RAM:clk, VGA_PLL:refclk, VGA_SUBSYSTEM:sys_clk_clk, VIDEO_DMA_ADDRESS_TRANSLATOR:clk, mm_interconnect_0:SYSTEM_PLL_sys_clk_clk, mm_interconnect_1:SYSTEM_PLL_sys_clk_clk, mm_interconnect_2:SYSTEM_PLL_sys_clk_clk, mm_interconnect_3:SYSTEM_PLL_sys_clk_clk, mm_interconnect_4:SYSTEM_PLL_sys_clk_clk, rst_controller:clk, rst_controller_003:clk]
	wire         dma_1_avalon_dma_master_waitrequest;                                // mm_interconnect_0:DMA_1_avalon_dma_master_waitrequest -> DMA_1:master_waitrequest
	wire   [7:0] dma_1_avalon_dma_master_readdata;                                   // mm_interconnect_0:DMA_1_avalon_dma_master_readdata -> DMA_1:master_readdata
	wire  [31:0] dma_1_avalon_dma_master_address;                                    // DMA_1:master_address -> mm_interconnect_0:DMA_1_avalon_dma_master_address
	wire         dma_1_avalon_dma_master_read;                                       // DMA_1:master_read -> mm_interconnect_0:DMA_1_avalon_dma_master_read
	wire         dma_1_avalon_dma_master_readdatavalid;                              // mm_interconnect_0:DMA_1_avalon_dma_master_readdatavalid -> DMA_1:master_readdatavalid
	wire         dma_1_avalon_dma_master_lock;                                       // DMA_1:master_arbiterlock -> mm_interconnect_0:DMA_1_avalon_dma_master_lock
	wire         dma_2_avalon_dma_master_waitrequest;                                // mm_interconnect_0:DMA_2_avalon_dma_master_waitrequest -> DMA_2:master_waitrequest
	wire   [7:0] dma_2_avalon_dma_master_readdata;                                   // mm_interconnect_0:DMA_2_avalon_dma_master_readdata -> DMA_2:master_readdata
	wire  [31:0] dma_2_avalon_dma_master_address;                                    // DMA_2:master_address -> mm_interconnect_0:DMA_2_avalon_dma_master_address
	wire         dma_2_avalon_dma_master_read;                                       // DMA_2:master_read -> mm_interconnect_0:DMA_2_avalon_dma_master_read
	wire         dma_2_avalon_dma_master_readdatavalid;                              // mm_interconnect_0:DMA_2_avalon_dma_master_readdatavalid -> DMA_2:master_readdatavalid
	wire         dma_2_avalon_dma_master_lock;                                       // DMA_2:master_arbiterlock -> mm_interconnect_0:DMA_2_avalon_dma_master_lock
	wire   [1:0] mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awburst;                 // mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_awburst -> ARM_A9_HPS:f2h_AWBURST
	wire   [4:0] mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awuser;                  // mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_awuser -> ARM_A9_HPS:f2h_AWUSER
	wire   [3:0] mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arlen;                   // mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_arlen -> ARM_A9_HPS:f2h_ARLEN
	wire   [7:0] mm_interconnect_0_arm_a9_hps_f2h_axi_slave_wstrb;                   // mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_wstrb -> ARM_A9_HPS:f2h_WSTRB
	wire         mm_interconnect_0_arm_a9_hps_f2h_axi_slave_wready;                  // ARM_A9_HPS:f2h_WREADY -> mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_wready
	wire   [7:0] mm_interconnect_0_arm_a9_hps_f2h_axi_slave_rid;                     // ARM_A9_HPS:f2h_RID -> mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_rid
	wire         mm_interconnect_0_arm_a9_hps_f2h_axi_slave_rready;                  // mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_rready -> ARM_A9_HPS:f2h_RREADY
	wire   [3:0] mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awlen;                   // mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_awlen -> ARM_A9_HPS:f2h_AWLEN
	wire   [7:0] mm_interconnect_0_arm_a9_hps_f2h_axi_slave_wid;                     // mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_wid -> ARM_A9_HPS:f2h_WID
	wire   [3:0] mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arcache;                 // mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_arcache -> ARM_A9_HPS:f2h_ARCACHE
	wire         mm_interconnect_0_arm_a9_hps_f2h_axi_slave_wvalid;                  // mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_wvalid -> ARM_A9_HPS:f2h_WVALID
	wire  [31:0] mm_interconnect_0_arm_a9_hps_f2h_axi_slave_araddr;                  // mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_araddr -> ARM_A9_HPS:f2h_ARADDR
	wire   [2:0] mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arprot;                  // mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_arprot -> ARM_A9_HPS:f2h_ARPROT
	wire   [2:0] mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awprot;                  // mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_awprot -> ARM_A9_HPS:f2h_AWPROT
	wire  [63:0] mm_interconnect_0_arm_a9_hps_f2h_axi_slave_wdata;                   // mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_wdata -> ARM_A9_HPS:f2h_WDATA
	wire         mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arvalid;                 // mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_arvalid -> ARM_A9_HPS:f2h_ARVALID
	wire   [3:0] mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awcache;                 // mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_awcache -> ARM_A9_HPS:f2h_AWCACHE
	wire   [7:0] mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arid;                    // mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_arid -> ARM_A9_HPS:f2h_ARID
	wire   [1:0] mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arlock;                  // mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_arlock -> ARM_A9_HPS:f2h_ARLOCK
	wire   [1:0] mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awlock;                  // mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_awlock -> ARM_A9_HPS:f2h_AWLOCK
	wire  [31:0] mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awaddr;                  // mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_awaddr -> ARM_A9_HPS:f2h_AWADDR
	wire   [1:0] mm_interconnect_0_arm_a9_hps_f2h_axi_slave_bresp;                   // ARM_A9_HPS:f2h_BRESP -> mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_bresp
	wire         mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arready;                 // ARM_A9_HPS:f2h_ARREADY -> mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_arready
	wire  [63:0] mm_interconnect_0_arm_a9_hps_f2h_axi_slave_rdata;                   // ARM_A9_HPS:f2h_RDATA -> mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_rdata
	wire         mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awready;                 // ARM_A9_HPS:f2h_AWREADY -> mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_awready
	wire   [1:0] mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arburst;                 // mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_arburst -> ARM_A9_HPS:f2h_ARBURST
	wire   [2:0] mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arsize;                  // mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_arsize -> ARM_A9_HPS:f2h_ARSIZE
	wire         mm_interconnect_0_arm_a9_hps_f2h_axi_slave_bready;                  // mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_bready -> ARM_A9_HPS:f2h_BREADY
	wire         mm_interconnect_0_arm_a9_hps_f2h_axi_slave_rlast;                   // ARM_A9_HPS:f2h_RLAST -> mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_rlast
	wire         mm_interconnect_0_arm_a9_hps_f2h_axi_slave_wlast;                   // mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_wlast -> ARM_A9_HPS:f2h_WLAST
	wire   [1:0] mm_interconnect_0_arm_a9_hps_f2h_axi_slave_rresp;                   // ARM_A9_HPS:f2h_RRESP -> mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_rresp
	wire   [7:0] mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awid;                    // mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_awid -> ARM_A9_HPS:f2h_AWID
	wire   [7:0] mm_interconnect_0_arm_a9_hps_f2h_axi_slave_bid;                     // ARM_A9_HPS:f2h_BID -> mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_bid
	wire         mm_interconnect_0_arm_a9_hps_f2h_axi_slave_bvalid;                  // ARM_A9_HPS:f2h_BVALID -> mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_bvalid
	wire   [2:0] mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awsize;                  // mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_awsize -> ARM_A9_HPS:f2h_AWSIZE
	wire         mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awvalid;                 // mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_awvalid -> ARM_A9_HPS:f2h_AWVALID
	wire   [4:0] mm_interconnect_0_arm_a9_hps_f2h_axi_slave_aruser;                  // mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_aruser -> ARM_A9_HPS:f2h_ARUSER
	wire         mm_interconnect_0_arm_a9_hps_f2h_axi_slave_rvalid;                  // ARM_A9_HPS:f2h_RVALID -> mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_rvalid
	wire         dma_write_avalon_dma_master_waitrequest;                            // mm_interconnect_1:DMA_WRITE_avalon_dma_master_waitrequest -> DMA_WRITE:master_waitrequest
	wire  [31:0] dma_write_avalon_dma_master_address;                                // DMA_WRITE:master_address -> mm_interconnect_1:DMA_WRITE_avalon_dma_master_address
	wire         dma_write_avalon_dma_master_write;                                  // DMA_WRITE:master_write -> mm_interconnect_1:DMA_WRITE_avalon_dma_master_write
	wire   [7:0] dma_write_avalon_dma_master_writedata;                              // DMA_WRITE:master_writedata -> mm_interconnect_1:DMA_WRITE_avalon_dma_master_writedata
	wire         mm_interconnect_1_ram_s1_chipselect;                                // mm_interconnect_1:RAM_s1_chipselect -> RAM:chipselect
	wire   [7:0] mm_interconnect_1_ram_s1_readdata;                                  // RAM:readdata -> mm_interconnect_1:RAM_s1_readdata
	wire  [18:0] mm_interconnect_1_ram_s1_address;                                   // mm_interconnect_1:RAM_s1_address -> RAM:address
	wire         mm_interconnect_1_ram_s1_write;                                     // mm_interconnect_1:RAM_s1_write -> RAM:write
	wire   [7:0] mm_interconnect_1_ram_s1_writedata;                                 // mm_interconnect_1:RAM_s1_writedata -> RAM:writedata
	wire         mm_interconnect_1_ram_s1_clken;                                     // mm_interconnect_1:RAM_s1_clken -> RAM:clken
	wire   [1:0] arm_a9_hps_h2f_lw_axi_master_awburst;                               // ARM_A9_HPS:h2f_lw_AWBURST -> mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_awburst
	wire   [3:0] arm_a9_hps_h2f_lw_axi_master_arlen;                                 // ARM_A9_HPS:h2f_lw_ARLEN -> mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_arlen
	wire   [3:0] arm_a9_hps_h2f_lw_axi_master_wstrb;                                 // ARM_A9_HPS:h2f_lw_WSTRB -> mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_wstrb
	wire         arm_a9_hps_h2f_lw_axi_master_wready;                                // mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_wready -> ARM_A9_HPS:h2f_lw_WREADY
	wire  [11:0] arm_a9_hps_h2f_lw_axi_master_rid;                                   // mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_rid -> ARM_A9_HPS:h2f_lw_RID
	wire         arm_a9_hps_h2f_lw_axi_master_rready;                                // ARM_A9_HPS:h2f_lw_RREADY -> mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_rready
	wire   [3:0] arm_a9_hps_h2f_lw_axi_master_awlen;                                 // ARM_A9_HPS:h2f_lw_AWLEN -> mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_awlen
	wire  [11:0] arm_a9_hps_h2f_lw_axi_master_wid;                                   // ARM_A9_HPS:h2f_lw_WID -> mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_wid
	wire   [3:0] arm_a9_hps_h2f_lw_axi_master_arcache;                               // ARM_A9_HPS:h2f_lw_ARCACHE -> mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_arcache
	wire         arm_a9_hps_h2f_lw_axi_master_wvalid;                                // ARM_A9_HPS:h2f_lw_WVALID -> mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_wvalid
	wire  [20:0] arm_a9_hps_h2f_lw_axi_master_araddr;                                // ARM_A9_HPS:h2f_lw_ARADDR -> mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_araddr
	wire   [2:0] arm_a9_hps_h2f_lw_axi_master_arprot;                                // ARM_A9_HPS:h2f_lw_ARPROT -> mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_arprot
	wire   [2:0] arm_a9_hps_h2f_lw_axi_master_awprot;                                // ARM_A9_HPS:h2f_lw_AWPROT -> mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_awprot
	wire  [31:0] arm_a9_hps_h2f_lw_axi_master_wdata;                                 // ARM_A9_HPS:h2f_lw_WDATA -> mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_wdata
	wire         arm_a9_hps_h2f_lw_axi_master_arvalid;                               // ARM_A9_HPS:h2f_lw_ARVALID -> mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_arvalid
	wire   [3:0] arm_a9_hps_h2f_lw_axi_master_awcache;                               // ARM_A9_HPS:h2f_lw_AWCACHE -> mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_awcache
	wire  [11:0] arm_a9_hps_h2f_lw_axi_master_arid;                                  // ARM_A9_HPS:h2f_lw_ARID -> mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_arid
	wire   [1:0] arm_a9_hps_h2f_lw_axi_master_arlock;                                // ARM_A9_HPS:h2f_lw_ARLOCK -> mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_arlock
	wire   [1:0] arm_a9_hps_h2f_lw_axi_master_awlock;                                // ARM_A9_HPS:h2f_lw_AWLOCK -> mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_awlock
	wire  [20:0] arm_a9_hps_h2f_lw_axi_master_awaddr;                                // ARM_A9_HPS:h2f_lw_AWADDR -> mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_awaddr
	wire   [1:0] arm_a9_hps_h2f_lw_axi_master_bresp;                                 // mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_bresp -> ARM_A9_HPS:h2f_lw_BRESP
	wire         arm_a9_hps_h2f_lw_axi_master_arready;                               // mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_arready -> ARM_A9_HPS:h2f_lw_ARREADY
	wire  [31:0] arm_a9_hps_h2f_lw_axi_master_rdata;                                 // mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_rdata -> ARM_A9_HPS:h2f_lw_RDATA
	wire         arm_a9_hps_h2f_lw_axi_master_awready;                               // mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_awready -> ARM_A9_HPS:h2f_lw_AWREADY
	wire   [1:0] arm_a9_hps_h2f_lw_axi_master_arburst;                               // ARM_A9_HPS:h2f_lw_ARBURST -> mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_arburst
	wire   [2:0] arm_a9_hps_h2f_lw_axi_master_arsize;                                // ARM_A9_HPS:h2f_lw_ARSIZE -> mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_arsize
	wire         arm_a9_hps_h2f_lw_axi_master_bready;                                // ARM_A9_HPS:h2f_lw_BREADY -> mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_bready
	wire         arm_a9_hps_h2f_lw_axi_master_rlast;                                 // mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_rlast -> ARM_A9_HPS:h2f_lw_RLAST
	wire         arm_a9_hps_h2f_lw_axi_master_wlast;                                 // ARM_A9_HPS:h2f_lw_WLAST -> mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_wlast
	wire   [1:0] arm_a9_hps_h2f_lw_axi_master_rresp;                                 // mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_rresp -> ARM_A9_HPS:h2f_lw_RRESP
	wire  [11:0] arm_a9_hps_h2f_lw_axi_master_awid;                                  // ARM_A9_HPS:h2f_lw_AWID -> mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_awid
	wire  [11:0] arm_a9_hps_h2f_lw_axi_master_bid;                                   // mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_bid -> ARM_A9_HPS:h2f_lw_BID
	wire         arm_a9_hps_h2f_lw_axi_master_bvalid;                                // mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_bvalid -> ARM_A9_HPS:h2f_lw_BVALID
	wire   [2:0] arm_a9_hps_h2f_lw_axi_master_awsize;                                // ARM_A9_HPS:h2f_lw_AWSIZE -> mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_awsize
	wire         arm_a9_hps_h2f_lw_axi_master_awvalid;                               // ARM_A9_HPS:h2f_lw_AWVALID -> mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_awvalid
	wire         arm_a9_hps_h2f_lw_axi_master_rvalid;                                // mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_rvalid -> ARM_A9_HPS:h2f_lw_RVALID
	wire  [31:0] mm_interconnect_2_dma_1_avalon_dma_control_slave_readdata;          // DMA_1:slave_readdata -> mm_interconnect_2:DMA_1_avalon_dma_control_slave_readdata
	wire   [1:0] mm_interconnect_2_dma_1_avalon_dma_control_slave_address;           // mm_interconnect_2:DMA_1_avalon_dma_control_slave_address -> DMA_1:slave_address
	wire         mm_interconnect_2_dma_1_avalon_dma_control_slave_read;              // mm_interconnect_2:DMA_1_avalon_dma_control_slave_read -> DMA_1:slave_read
	wire   [3:0] mm_interconnect_2_dma_1_avalon_dma_control_slave_byteenable;        // mm_interconnect_2:DMA_1_avalon_dma_control_slave_byteenable -> DMA_1:slave_byteenable
	wire         mm_interconnect_2_dma_1_avalon_dma_control_slave_write;             // mm_interconnect_2:DMA_1_avalon_dma_control_slave_write -> DMA_1:slave_write
	wire  [31:0] mm_interconnect_2_dma_1_avalon_dma_control_slave_writedata;         // mm_interconnect_2:DMA_1_avalon_dma_control_slave_writedata -> DMA_1:slave_writedata
	wire  [31:0] mm_interconnect_2_dma_2_avalon_dma_control_slave_readdata;          // DMA_2:slave_readdata -> mm_interconnect_2:DMA_2_avalon_dma_control_slave_readdata
	wire   [1:0] mm_interconnect_2_dma_2_avalon_dma_control_slave_address;           // mm_interconnect_2:DMA_2_avalon_dma_control_slave_address -> DMA_2:slave_address
	wire         mm_interconnect_2_dma_2_avalon_dma_control_slave_read;              // mm_interconnect_2:DMA_2_avalon_dma_control_slave_read -> DMA_2:slave_read
	wire   [3:0] mm_interconnect_2_dma_2_avalon_dma_control_slave_byteenable;        // mm_interconnect_2:DMA_2_avalon_dma_control_slave_byteenable -> DMA_2:slave_byteenable
	wire         mm_interconnect_2_dma_2_avalon_dma_control_slave_write;             // mm_interconnect_2:DMA_2_avalon_dma_control_slave_write -> DMA_2:slave_write
	wire  [31:0] mm_interconnect_2_dma_2_avalon_dma_control_slave_writedata;         // mm_interconnect_2:DMA_2_avalon_dma_control_slave_writedata -> DMA_2:slave_writedata
	wire  [31:0] mm_interconnect_2_dma_write_avalon_dma_control_slave_readdata;      // DMA_WRITE:slave_readdata -> mm_interconnect_2:DMA_WRITE_avalon_dma_control_slave_readdata
	wire   [1:0] mm_interconnect_2_dma_write_avalon_dma_control_slave_address;       // mm_interconnect_2:DMA_WRITE_avalon_dma_control_slave_address -> DMA_WRITE:slave_address
	wire         mm_interconnect_2_dma_write_avalon_dma_control_slave_read;          // mm_interconnect_2:DMA_WRITE_avalon_dma_control_slave_read -> DMA_WRITE:slave_read
	wire   [3:0] mm_interconnect_2_dma_write_avalon_dma_control_slave_byteenable;    // mm_interconnect_2:DMA_WRITE_avalon_dma_control_slave_byteenable -> DMA_WRITE:slave_byteenable
	wire         mm_interconnect_2_dma_write_avalon_dma_control_slave_write;         // mm_interconnect_2:DMA_WRITE_avalon_dma_control_slave_write -> DMA_WRITE:slave_write
	wire  [31:0] mm_interconnect_2_dma_write_avalon_dma_control_slave_writedata;     // mm_interconnect_2:DMA_WRITE_avalon_dma_control_slave_writedata -> DMA_WRITE:slave_writedata
	wire  [31:0] mm_interconnect_2_video_dma_address_translator_slave_readdata;      // VIDEO_DMA_ADDRESS_TRANSLATOR:slave_readdata -> mm_interconnect_2:VIDEO_DMA_ADDRESS_TRANSLATOR_slave_readdata
	wire         mm_interconnect_2_video_dma_address_translator_slave_waitrequest;   // VIDEO_DMA_ADDRESS_TRANSLATOR:slave_waitrequest -> mm_interconnect_2:VIDEO_DMA_ADDRESS_TRANSLATOR_slave_waitrequest
	wire   [1:0] mm_interconnect_2_video_dma_address_translator_slave_address;       // mm_interconnect_2:VIDEO_DMA_ADDRESS_TRANSLATOR_slave_address -> VIDEO_DMA_ADDRESS_TRANSLATOR:slave_address
	wire         mm_interconnect_2_video_dma_address_translator_slave_read;          // mm_interconnect_2:VIDEO_DMA_ADDRESS_TRANSLATOR_slave_read -> VIDEO_DMA_ADDRESS_TRANSLATOR:slave_read
	wire   [3:0] mm_interconnect_2_video_dma_address_translator_slave_byteenable;    // mm_interconnect_2:VIDEO_DMA_ADDRESS_TRANSLATOR_slave_byteenable -> VIDEO_DMA_ADDRESS_TRANSLATOR:slave_byteenable
	wire         mm_interconnect_2_video_dma_address_translator_slave_write;         // mm_interconnect_2:VIDEO_DMA_ADDRESS_TRANSLATOR_slave_write -> VIDEO_DMA_ADDRESS_TRANSLATOR:slave_write
	wire  [31:0] mm_interconnect_2_video_dma_address_translator_slave_writedata;     // mm_interconnect_2:VIDEO_DMA_ADDRESS_TRANSLATOR_slave_writedata -> VIDEO_DMA_ADDRESS_TRANSLATOR:slave_writedata
	wire  [31:0] video_dma_address_translator_master_readdata;                       // mm_interconnect_3:VIDEO_DMA_ADDRESS_TRANSLATOR_master_readdata -> VIDEO_DMA_ADDRESS_TRANSLATOR:master_readdata
	wire         video_dma_address_translator_master_waitrequest;                    // mm_interconnect_3:VIDEO_DMA_ADDRESS_TRANSLATOR_master_waitrequest -> VIDEO_DMA_ADDRESS_TRANSLATOR:master_waitrequest
	wire   [1:0] video_dma_address_translator_master_address;                        // VIDEO_DMA_ADDRESS_TRANSLATOR:master_address -> mm_interconnect_3:VIDEO_DMA_ADDRESS_TRANSLATOR_master_address
	wire   [3:0] video_dma_address_translator_master_byteenable;                     // VIDEO_DMA_ADDRESS_TRANSLATOR:master_byteenable -> mm_interconnect_3:VIDEO_DMA_ADDRESS_TRANSLATOR_master_byteenable
	wire         video_dma_address_translator_master_read;                           // VIDEO_DMA_ADDRESS_TRANSLATOR:master_read -> mm_interconnect_3:VIDEO_DMA_ADDRESS_TRANSLATOR_master_read
	wire         video_dma_address_translator_master_write;                          // VIDEO_DMA_ADDRESS_TRANSLATOR:master_write -> mm_interconnect_3:VIDEO_DMA_ADDRESS_TRANSLATOR_master_write
	wire  [31:0] video_dma_address_translator_master_writedata;                      // VIDEO_DMA_ADDRESS_TRANSLATOR:master_writedata -> mm_interconnect_3:VIDEO_DMA_ADDRESS_TRANSLATOR_master_writedata
	wire  [31:0] mm_interconnect_3_vga_subsystem_pixel_dma_control_slave_readdata;   // VGA_SUBSYSTEM:pixel_dma_control_slave_readdata -> mm_interconnect_3:VGA_SUBSYSTEM_pixel_dma_control_slave_readdata
	wire   [1:0] mm_interconnect_3_vga_subsystem_pixel_dma_control_slave_address;    // mm_interconnect_3:VGA_SUBSYSTEM_pixel_dma_control_slave_address -> VGA_SUBSYSTEM:pixel_dma_control_slave_address
	wire         mm_interconnect_3_vga_subsystem_pixel_dma_control_slave_read;       // mm_interconnect_3:VGA_SUBSYSTEM_pixel_dma_control_slave_read -> VGA_SUBSYSTEM:pixel_dma_control_slave_read
	wire   [3:0] mm_interconnect_3_vga_subsystem_pixel_dma_control_slave_byteenable; // mm_interconnect_3:VGA_SUBSYSTEM_pixel_dma_control_slave_byteenable -> VGA_SUBSYSTEM:pixel_dma_control_slave_byteenable
	wire         mm_interconnect_3_vga_subsystem_pixel_dma_control_slave_write;      // mm_interconnect_3:VGA_SUBSYSTEM_pixel_dma_control_slave_write -> VGA_SUBSYSTEM:pixel_dma_control_slave_write
	wire  [31:0] mm_interconnect_3_vga_subsystem_pixel_dma_control_slave_writedata;  // mm_interconnect_3:VGA_SUBSYSTEM_pixel_dma_control_slave_writedata -> VGA_SUBSYSTEM:pixel_dma_control_slave_writedata
	wire         vga_subsystem_pixel_dma_master_waitrequest;                         // mm_interconnect_4:VGA_SUBSYSTEM_pixel_dma_master_waitrequest -> VGA_SUBSYSTEM:pixel_dma_master_waitrequest
	wire   [7:0] vga_subsystem_pixel_dma_master_readdata;                            // mm_interconnect_4:VGA_SUBSYSTEM_pixel_dma_master_readdata -> VGA_SUBSYSTEM:pixel_dma_master_readdata
	wire  [31:0] vga_subsystem_pixel_dma_master_address;                             // VGA_SUBSYSTEM:pixel_dma_master_address -> mm_interconnect_4:VGA_SUBSYSTEM_pixel_dma_master_address
	wire         vga_subsystem_pixel_dma_master_read;                                // VGA_SUBSYSTEM:pixel_dma_master_read -> mm_interconnect_4:VGA_SUBSYSTEM_pixel_dma_master_read
	wire         vga_subsystem_pixel_dma_master_readdatavalid;                       // mm_interconnect_4:VGA_SUBSYSTEM_pixel_dma_master_readdatavalid -> VGA_SUBSYSTEM:pixel_dma_master_readdatavalid
	wire         vga_subsystem_pixel_dma_master_lock;                                // VGA_SUBSYSTEM:pixel_dma_master_lock -> mm_interconnect_4:VGA_SUBSYSTEM_pixel_dma_master_lock
	wire         mm_interconnect_4_ram_s2_chipselect;                                // mm_interconnect_4:RAM_s2_chipselect -> RAM:chipselect2
	wire   [7:0] mm_interconnect_4_ram_s2_readdata;                                  // RAM:readdata2 -> mm_interconnect_4:RAM_s2_readdata
	wire  [18:0] mm_interconnect_4_ram_s2_address;                                   // mm_interconnect_4:RAM_s2_address -> RAM:address2
	wire         mm_interconnect_4_ram_s2_write;                                     // mm_interconnect_4:RAM_s2_write -> RAM:write2
	wire   [7:0] mm_interconnect_4_ram_s2_writedata;                                 // mm_interconnect_4:RAM_s2_writedata -> RAM:writedata2
	wire         mm_interconnect_4_ram_s2_clken;                                     // mm_interconnect_4:RAM_s2_clken -> RAM:clken2
	wire  [31:0] arm_a9_hps_f2h_irq0_irq;                                            // irq_mapper:sender_irq -> ARM_A9_HPS:f2h_irq_p0
	wire  [31:0] arm_a9_hps_f2h_irq1_irq;                                            // irq_mapper_001:sender_irq -> ARM_A9_HPS:f2h_irq_p1
	wire         rst_controller_reset_out_reset;                                     // rst_controller:reset_out -> [BUFFER_1:reset, BUFFER_2:reset, DMA_1:reset, DMA_2:reset, DMA_WRITE:reset, FUSION:reset, PADDING_1:reset, PADDING_2:reset, RAM:reset, VIDEO_DMA_ADDRESS_TRANSLATOR:reset, mm_interconnect_0:DMA_1_reset_reset_bridge_in_reset_reset, mm_interconnect_1:DMA_WRITE_reset_reset_bridge_in_reset_reset, mm_interconnect_2:DMA_1_reset_reset_bridge_in_reset_reset, mm_interconnect_3:VGA_SUBSYSTEM_sys_reset_reset_bridge_in_reset_reset, mm_interconnect_3:VIDEO_DMA_ADDRESS_TRANSLATOR_reset_reset_bridge_in_reset_reset, mm_interconnect_4:RAM_reset1_reset_bridge_in_reset_reset, mm_interconnect_4:VGA_SUBSYSTEM_sys_reset_reset_bridge_in_reset_reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                                 // rst_controller:reset_req -> [RAM:reset_req, rst_translator:reset_req_in]
	wire         arm_a9_hps_h2f_reset_reset;                                         // ARM_A9_HPS:h2f_rst_n -> [rst_controller:reset_in0, rst_controller_001:reset_in0, rst_controller_002:reset_in0, rst_controller_003:reset_in0]
	wire         system_pll_reset_source_reset;                                      // SYSTEM_PLL:reset_source_reset -> [rst_controller:reset_in1, rst_controller_001:reset_in1, rst_controller_002:reset_in1]
	wire         rst_controller_001_reset_out_reset;                                 // rst_controller_001:reset_out -> VGA_PLL:rst
	wire         rst_controller_002_reset_out_reset;                                 // rst_controller_002:reset_out -> VGA_SUBSYSTEM:sys_reset_reset_n
	wire         rst_controller_003_reset_out_reset;                                 // rst_controller_003:reset_out -> [mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset]

	Computer_System_ARM_A9_HPS #(
		.F2S_Width (2),
		.S2F_Width (3)
	) arm_a9_hps (
		.mem_a                    (memory_mem_a),                                       //            memory.mem_a
		.mem_ba                   (memory_mem_ba),                                      //                  .mem_ba
		.mem_ck                   (memory_mem_ck),                                      //                  .mem_ck
		.mem_ck_n                 (memory_mem_ck_n),                                    //                  .mem_ck_n
		.mem_cke                  (memory_mem_cke),                                     //                  .mem_cke
		.mem_cs_n                 (memory_mem_cs_n),                                    //                  .mem_cs_n
		.mem_ras_n                (memory_mem_ras_n),                                   //                  .mem_ras_n
		.mem_cas_n                (memory_mem_cas_n),                                   //                  .mem_cas_n
		.mem_we_n                 (memory_mem_we_n),                                    //                  .mem_we_n
		.mem_reset_n              (memory_mem_reset_n),                                 //                  .mem_reset_n
		.mem_dq                   (memory_mem_dq),                                      //                  .mem_dq
		.mem_dqs                  (memory_mem_dqs),                                     //                  .mem_dqs
		.mem_dqs_n                (memory_mem_dqs_n),                                   //                  .mem_dqs_n
		.mem_odt                  (memory_mem_odt),                                     //                  .mem_odt
		.mem_dm                   (memory_mem_dm),                                      //                  .mem_dm
		.oct_rzqin                (memory_oct_rzqin),                                   //                  .oct_rzqin
		.hps_io_emac1_inst_TX_CLK (hps_io_hps_io_emac1_inst_TX_CLK),                    //            hps_io.hps_io_emac1_inst_TX_CLK
		.hps_io_emac1_inst_TXD0   (hps_io_hps_io_emac1_inst_TXD0),                      //                  .hps_io_emac1_inst_TXD0
		.hps_io_emac1_inst_TXD1   (hps_io_hps_io_emac1_inst_TXD1),                      //                  .hps_io_emac1_inst_TXD1
		.hps_io_emac1_inst_TXD2   (hps_io_hps_io_emac1_inst_TXD2),                      //                  .hps_io_emac1_inst_TXD2
		.hps_io_emac1_inst_TXD3   (hps_io_hps_io_emac1_inst_TXD3),                      //                  .hps_io_emac1_inst_TXD3
		.hps_io_emac1_inst_RXD0   (hps_io_hps_io_emac1_inst_RXD0),                      //                  .hps_io_emac1_inst_RXD0
		.hps_io_emac1_inst_MDIO   (hps_io_hps_io_emac1_inst_MDIO),                      //                  .hps_io_emac1_inst_MDIO
		.hps_io_emac1_inst_MDC    (hps_io_hps_io_emac1_inst_MDC),                       //                  .hps_io_emac1_inst_MDC
		.hps_io_emac1_inst_RX_CTL (hps_io_hps_io_emac1_inst_RX_CTL),                    //                  .hps_io_emac1_inst_RX_CTL
		.hps_io_emac1_inst_TX_CTL (hps_io_hps_io_emac1_inst_TX_CTL),                    //                  .hps_io_emac1_inst_TX_CTL
		.hps_io_emac1_inst_RX_CLK (hps_io_hps_io_emac1_inst_RX_CLK),                    //                  .hps_io_emac1_inst_RX_CLK
		.hps_io_emac1_inst_RXD1   (hps_io_hps_io_emac1_inst_RXD1),                      //                  .hps_io_emac1_inst_RXD1
		.hps_io_emac1_inst_RXD2   (hps_io_hps_io_emac1_inst_RXD2),                      //                  .hps_io_emac1_inst_RXD2
		.hps_io_emac1_inst_RXD3   (hps_io_hps_io_emac1_inst_RXD3),                      //                  .hps_io_emac1_inst_RXD3
		.hps_io_qspi_inst_IO0     (hps_io_hps_io_qspi_inst_IO0),                        //                  .hps_io_qspi_inst_IO0
		.hps_io_qspi_inst_IO1     (hps_io_hps_io_qspi_inst_IO1),                        //                  .hps_io_qspi_inst_IO1
		.hps_io_qspi_inst_IO2     (hps_io_hps_io_qspi_inst_IO2),                        //                  .hps_io_qspi_inst_IO2
		.hps_io_qspi_inst_IO3     (hps_io_hps_io_qspi_inst_IO3),                        //                  .hps_io_qspi_inst_IO3
		.hps_io_qspi_inst_SS0     (hps_io_hps_io_qspi_inst_SS0),                        //                  .hps_io_qspi_inst_SS0
		.hps_io_qspi_inst_CLK     (hps_io_hps_io_qspi_inst_CLK),                        //                  .hps_io_qspi_inst_CLK
		.hps_io_sdio_inst_CMD     (hps_io_hps_io_sdio_inst_CMD),                        //                  .hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0      (hps_io_hps_io_sdio_inst_D0),                         //                  .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1      (hps_io_hps_io_sdio_inst_D1),                         //                  .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK     (hps_io_hps_io_sdio_inst_CLK),                        //                  .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2      (hps_io_hps_io_sdio_inst_D2),                         //                  .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3      (hps_io_hps_io_sdio_inst_D3),                         //                  .hps_io_sdio_inst_D3
		.hps_io_usb1_inst_D0      (hps_io_hps_io_usb1_inst_D0),                         //                  .hps_io_usb1_inst_D0
		.hps_io_usb1_inst_D1      (hps_io_hps_io_usb1_inst_D1),                         //                  .hps_io_usb1_inst_D1
		.hps_io_usb1_inst_D2      (hps_io_hps_io_usb1_inst_D2),                         //                  .hps_io_usb1_inst_D2
		.hps_io_usb1_inst_D3      (hps_io_hps_io_usb1_inst_D3),                         //                  .hps_io_usb1_inst_D3
		.hps_io_usb1_inst_D4      (hps_io_hps_io_usb1_inst_D4),                         //                  .hps_io_usb1_inst_D4
		.hps_io_usb1_inst_D5      (hps_io_hps_io_usb1_inst_D5),                         //                  .hps_io_usb1_inst_D5
		.hps_io_usb1_inst_D6      (hps_io_hps_io_usb1_inst_D6),                         //                  .hps_io_usb1_inst_D6
		.hps_io_usb1_inst_D7      (hps_io_hps_io_usb1_inst_D7),                         //                  .hps_io_usb1_inst_D7
		.hps_io_usb1_inst_CLK     (hps_io_hps_io_usb1_inst_CLK),                        //                  .hps_io_usb1_inst_CLK
		.hps_io_usb1_inst_STP     (hps_io_hps_io_usb1_inst_STP),                        //                  .hps_io_usb1_inst_STP
		.hps_io_usb1_inst_DIR     (hps_io_hps_io_usb1_inst_DIR),                        //                  .hps_io_usb1_inst_DIR
		.hps_io_usb1_inst_NXT     (hps_io_hps_io_usb1_inst_NXT),                        //                  .hps_io_usb1_inst_NXT
		.hps_io_spim1_inst_CLK    (hps_io_hps_io_spim1_inst_CLK),                       //                  .hps_io_spim1_inst_CLK
		.hps_io_spim1_inst_MOSI   (hps_io_hps_io_spim1_inst_MOSI),                      //                  .hps_io_spim1_inst_MOSI
		.hps_io_spim1_inst_MISO   (hps_io_hps_io_spim1_inst_MISO),                      //                  .hps_io_spim1_inst_MISO
		.hps_io_spim1_inst_SS0    (hps_io_hps_io_spim1_inst_SS0),                       //                  .hps_io_spim1_inst_SS0
		.hps_io_uart0_inst_RX     (hps_io_hps_io_uart0_inst_RX),                        //                  .hps_io_uart0_inst_RX
		.hps_io_uart0_inst_TX     (hps_io_hps_io_uart0_inst_TX),                        //                  .hps_io_uart0_inst_TX
		.hps_io_i2c0_inst_SDA     (hps_io_hps_io_i2c0_inst_SDA),                        //                  .hps_io_i2c0_inst_SDA
		.hps_io_i2c0_inst_SCL     (hps_io_hps_io_i2c0_inst_SCL),                        //                  .hps_io_i2c0_inst_SCL
		.hps_io_i2c1_inst_SDA     (hps_io_hps_io_i2c1_inst_SDA),                        //                  .hps_io_i2c1_inst_SDA
		.hps_io_i2c1_inst_SCL     (hps_io_hps_io_i2c1_inst_SCL),                        //                  .hps_io_i2c1_inst_SCL
		.hps_io_gpio_inst_GPIO09  (hps_io_hps_io_gpio_inst_GPIO09),                     //                  .hps_io_gpio_inst_GPIO09
		.hps_io_gpio_inst_GPIO35  (hps_io_hps_io_gpio_inst_GPIO35),                     //                  .hps_io_gpio_inst_GPIO35
		.hps_io_gpio_inst_GPIO40  (hps_io_hps_io_gpio_inst_GPIO40),                     //                  .hps_io_gpio_inst_GPIO40
		.hps_io_gpio_inst_GPIO41  (hps_io_hps_io_gpio_inst_GPIO41),                     //                  .hps_io_gpio_inst_GPIO41
		.hps_io_gpio_inst_GPIO48  (hps_io_hps_io_gpio_inst_GPIO48),                     //                  .hps_io_gpio_inst_GPIO48
		.hps_io_gpio_inst_GPIO53  (hps_io_hps_io_gpio_inst_GPIO53),                     //                  .hps_io_gpio_inst_GPIO53
		.hps_io_gpio_inst_GPIO54  (hps_io_hps_io_gpio_inst_GPIO54),                     //                  .hps_io_gpio_inst_GPIO54
		.hps_io_gpio_inst_GPIO61  (hps_io_hps_io_gpio_inst_GPIO61),                     //                  .hps_io_gpio_inst_GPIO61
		.h2f_rst_n                (arm_a9_hps_h2f_reset_reset),                         //         h2f_reset.reset_n
		.h2f_axi_clk              (system_pll_sys_clk_clk),                             //     h2f_axi_clock.clk
		.h2f_AWID                 (),                                                   //    h2f_axi_master.awid
		.h2f_AWADDR               (),                                                   //                  .awaddr
		.h2f_AWLEN                (),                                                   //                  .awlen
		.h2f_AWSIZE               (),                                                   //                  .awsize
		.h2f_AWBURST              (),                                                   //                  .awburst
		.h2f_AWLOCK               (),                                                   //                  .awlock
		.h2f_AWCACHE              (),                                                   //                  .awcache
		.h2f_AWPROT               (),                                                   //                  .awprot
		.h2f_AWVALID              (),                                                   //                  .awvalid
		.h2f_AWREADY              (),                                                   //                  .awready
		.h2f_WID                  (),                                                   //                  .wid
		.h2f_WDATA                (),                                                   //                  .wdata
		.h2f_WSTRB                (),                                                   //                  .wstrb
		.h2f_WLAST                (),                                                   //                  .wlast
		.h2f_WVALID               (),                                                   //                  .wvalid
		.h2f_WREADY               (),                                                   //                  .wready
		.h2f_BID                  (),                                                   //                  .bid
		.h2f_BRESP                (),                                                   //                  .bresp
		.h2f_BVALID               (),                                                   //                  .bvalid
		.h2f_BREADY               (),                                                   //                  .bready
		.h2f_ARID                 (),                                                   //                  .arid
		.h2f_ARADDR               (),                                                   //                  .araddr
		.h2f_ARLEN                (),                                                   //                  .arlen
		.h2f_ARSIZE               (),                                                   //                  .arsize
		.h2f_ARBURST              (),                                                   //                  .arburst
		.h2f_ARLOCK               (),                                                   //                  .arlock
		.h2f_ARCACHE              (),                                                   //                  .arcache
		.h2f_ARPROT               (),                                                   //                  .arprot
		.h2f_ARVALID              (),                                                   //                  .arvalid
		.h2f_ARREADY              (),                                                   //                  .arready
		.h2f_RID                  (),                                                   //                  .rid
		.h2f_RDATA                (),                                                   //                  .rdata
		.h2f_RRESP                (),                                                   //                  .rresp
		.h2f_RLAST                (),                                                   //                  .rlast
		.h2f_RVALID               (),                                                   //                  .rvalid
		.h2f_RREADY               (),                                                   //                  .rready
		.f2h_axi_clk              (system_pll_sys_clk_clk),                             //     f2h_axi_clock.clk
		.f2h_AWID                 (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awid),    //     f2h_axi_slave.awid
		.f2h_AWADDR               (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awaddr),  //                  .awaddr
		.f2h_AWLEN                (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awlen),   //                  .awlen
		.f2h_AWSIZE               (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awsize),  //                  .awsize
		.f2h_AWBURST              (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awburst), //                  .awburst
		.f2h_AWLOCK               (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awlock),  //                  .awlock
		.f2h_AWCACHE              (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awcache), //                  .awcache
		.f2h_AWPROT               (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awprot),  //                  .awprot
		.f2h_AWVALID              (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awvalid), //                  .awvalid
		.f2h_AWREADY              (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awready), //                  .awready
		.f2h_AWUSER               (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awuser),  //                  .awuser
		.f2h_WID                  (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_wid),     //                  .wid
		.f2h_WDATA                (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_wdata),   //                  .wdata
		.f2h_WSTRB                (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_wstrb),   //                  .wstrb
		.f2h_WLAST                (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_wlast),   //                  .wlast
		.f2h_WVALID               (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_wvalid),  //                  .wvalid
		.f2h_WREADY               (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_wready),  //                  .wready
		.f2h_BID                  (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_bid),     //                  .bid
		.f2h_BRESP                (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_bresp),   //                  .bresp
		.f2h_BVALID               (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_bvalid),  //                  .bvalid
		.f2h_BREADY               (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_bready),  //                  .bready
		.f2h_ARID                 (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arid),    //                  .arid
		.f2h_ARADDR               (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_araddr),  //                  .araddr
		.f2h_ARLEN                (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arlen),   //                  .arlen
		.f2h_ARSIZE               (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arsize),  //                  .arsize
		.f2h_ARBURST              (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arburst), //                  .arburst
		.f2h_ARLOCK               (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arlock),  //                  .arlock
		.f2h_ARCACHE              (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arcache), //                  .arcache
		.f2h_ARPROT               (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arprot),  //                  .arprot
		.f2h_ARVALID              (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arvalid), //                  .arvalid
		.f2h_ARREADY              (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arready), //                  .arready
		.f2h_ARUSER               (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_aruser),  //                  .aruser
		.f2h_RID                  (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_rid),     //                  .rid
		.f2h_RDATA                (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_rdata),   //                  .rdata
		.f2h_RRESP                (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_rresp),   //                  .rresp
		.f2h_RLAST                (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_rlast),   //                  .rlast
		.f2h_RVALID               (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_rvalid),  //                  .rvalid
		.f2h_RREADY               (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_rready),  //                  .rready
		.h2f_lw_axi_clk           (system_pll_sys_clk_clk),                             //  h2f_lw_axi_clock.clk
		.h2f_lw_AWID              (arm_a9_hps_h2f_lw_axi_master_awid),                  // h2f_lw_axi_master.awid
		.h2f_lw_AWADDR            (arm_a9_hps_h2f_lw_axi_master_awaddr),                //                  .awaddr
		.h2f_lw_AWLEN             (arm_a9_hps_h2f_lw_axi_master_awlen),                 //                  .awlen
		.h2f_lw_AWSIZE            (arm_a9_hps_h2f_lw_axi_master_awsize),                //                  .awsize
		.h2f_lw_AWBURST           (arm_a9_hps_h2f_lw_axi_master_awburst),               //                  .awburst
		.h2f_lw_AWLOCK            (arm_a9_hps_h2f_lw_axi_master_awlock),                //                  .awlock
		.h2f_lw_AWCACHE           (arm_a9_hps_h2f_lw_axi_master_awcache),               //                  .awcache
		.h2f_lw_AWPROT            (arm_a9_hps_h2f_lw_axi_master_awprot),                //                  .awprot
		.h2f_lw_AWVALID           (arm_a9_hps_h2f_lw_axi_master_awvalid),               //                  .awvalid
		.h2f_lw_AWREADY           (arm_a9_hps_h2f_lw_axi_master_awready),               //                  .awready
		.h2f_lw_WID               (arm_a9_hps_h2f_lw_axi_master_wid),                   //                  .wid
		.h2f_lw_WDATA             (arm_a9_hps_h2f_lw_axi_master_wdata),                 //                  .wdata
		.h2f_lw_WSTRB             (arm_a9_hps_h2f_lw_axi_master_wstrb),                 //                  .wstrb
		.h2f_lw_WLAST             (arm_a9_hps_h2f_lw_axi_master_wlast),                 //                  .wlast
		.h2f_lw_WVALID            (arm_a9_hps_h2f_lw_axi_master_wvalid),                //                  .wvalid
		.h2f_lw_WREADY            (arm_a9_hps_h2f_lw_axi_master_wready),                //                  .wready
		.h2f_lw_BID               (arm_a9_hps_h2f_lw_axi_master_bid),                   //                  .bid
		.h2f_lw_BRESP             (arm_a9_hps_h2f_lw_axi_master_bresp),                 //                  .bresp
		.h2f_lw_BVALID            (arm_a9_hps_h2f_lw_axi_master_bvalid),                //                  .bvalid
		.h2f_lw_BREADY            (arm_a9_hps_h2f_lw_axi_master_bready),                //                  .bready
		.h2f_lw_ARID              (arm_a9_hps_h2f_lw_axi_master_arid),                  //                  .arid
		.h2f_lw_ARADDR            (arm_a9_hps_h2f_lw_axi_master_araddr),                //                  .araddr
		.h2f_lw_ARLEN             (arm_a9_hps_h2f_lw_axi_master_arlen),                 //                  .arlen
		.h2f_lw_ARSIZE            (arm_a9_hps_h2f_lw_axi_master_arsize),                //                  .arsize
		.h2f_lw_ARBURST           (arm_a9_hps_h2f_lw_axi_master_arburst),               //                  .arburst
		.h2f_lw_ARLOCK            (arm_a9_hps_h2f_lw_axi_master_arlock),                //                  .arlock
		.h2f_lw_ARCACHE           (arm_a9_hps_h2f_lw_axi_master_arcache),               //                  .arcache
		.h2f_lw_ARPROT            (arm_a9_hps_h2f_lw_axi_master_arprot),                //                  .arprot
		.h2f_lw_ARVALID           (arm_a9_hps_h2f_lw_axi_master_arvalid),               //                  .arvalid
		.h2f_lw_ARREADY           (arm_a9_hps_h2f_lw_axi_master_arready),               //                  .arready
		.h2f_lw_RID               (arm_a9_hps_h2f_lw_axi_master_rid),                   //                  .rid
		.h2f_lw_RDATA             (arm_a9_hps_h2f_lw_axi_master_rdata),                 //                  .rdata
		.h2f_lw_RRESP             (arm_a9_hps_h2f_lw_axi_master_rresp),                 //                  .rresp
		.h2f_lw_RLAST             (arm_a9_hps_h2f_lw_axi_master_rlast),                 //                  .rlast
		.h2f_lw_RVALID            (arm_a9_hps_h2f_lw_axi_master_rvalid),                //                  .rvalid
		.h2f_lw_RREADY            (arm_a9_hps_h2f_lw_axi_master_rready),                //                  .rready
		.f2h_irq_p0               (arm_a9_hps_f2h_irq0_irq),                            //          f2h_irq0.irq
		.f2h_irq_p1               (arm_a9_hps_f2h_irq1_irq)                             //          f2h_irq1.irq
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (8),
		.FIFO_DEPTH          (8192),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (3),
		.USE_MEMORY_BLOCKS   (1),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) buffer_1 (
		.clk               (system_pll_sys_clk_clk),                  //       clk.clk
		.reset             (rst_controller_reset_out_reset),          // clk_reset.reset
		.in_data           (dma_1_avalon_pixel_source_data),          //        in.data
		.in_valid          (dma_1_avalon_pixel_source_valid),         //          .valid
		.in_ready          (dma_1_avalon_pixel_source_ready),         //          .ready
		.in_startofpacket  (dma_1_avalon_pixel_source_startofpacket), //          .startofpacket
		.in_endofpacket    (dma_1_avalon_pixel_source_endofpacket),   //          .endofpacket
		.out_data          (buffer_1_out_data),                       //       out.data
		.out_valid         (buffer_1_out_valid),                      //          .valid
		.out_ready         (buffer_1_out_ready),                      //          .ready
		.out_startofpacket (buffer_1_out_startofpacket),              //          .startofpacket
		.out_endofpacket   (buffer_1_out_endofpacket),                //          .endofpacket
		.csr_address       (2'b00),                                   // (terminated)
		.csr_read          (1'b0),                                    // (terminated)
		.csr_write         (1'b0),                                    // (terminated)
		.csr_readdata      (),                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),    // (terminated)
		.almost_full_data  (),                                        // (terminated)
		.almost_empty_data (),                                        // (terminated)
		.in_empty          (1'b0),                                    // (terminated)
		.out_empty         (),                                        // (terminated)
		.in_error          (1'b0),                                    // (terminated)
		.out_error         (),                                        // (terminated)
		.in_channel        (1'b0),                                    // (terminated)
		.out_channel       ()                                         // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (8),
		.FIFO_DEPTH          (8192),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (3),
		.USE_MEMORY_BLOCKS   (1),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) buffer_2 (
		.clk               (system_pll_sys_clk_clk),                  //       clk.clk
		.reset             (rst_controller_reset_out_reset),          // clk_reset.reset
		.in_data           (dma_2_avalon_pixel_source_data),          //        in.data
		.in_valid          (dma_2_avalon_pixel_source_valid),         //          .valid
		.in_ready          (dma_2_avalon_pixel_source_ready),         //          .ready
		.in_startofpacket  (dma_2_avalon_pixel_source_startofpacket), //          .startofpacket
		.in_endofpacket    (dma_2_avalon_pixel_source_endofpacket),   //          .endofpacket
		.out_data          (buffer_2_out_data),                       //       out.data
		.out_valid         (buffer_2_out_valid),                      //          .valid
		.out_ready         (buffer_2_out_ready),                      //          .ready
		.out_startofpacket (buffer_2_out_startofpacket),              //          .startofpacket
		.out_endofpacket   (buffer_2_out_endofpacket),                //          .endofpacket
		.csr_address       (2'b00),                                   // (terminated)
		.csr_read          (1'b0),                                    // (terminated)
		.csr_write         (1'b0),                                    // (terminated)
		.csr_readdata      (),                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),    // (terminated)
		.almost_full_data  (),                                        // (terminated)
		.almost_empty_data (),                                        // (terminated)
		.in_empty          (1'b0),                                    // (terminated)
		.out_empty         (),                                        // (terminated)
		.in_error          (1'b0),                                    // (terminated)
		.out_error         (),                                        // (terminated)
		.in_channel        (1'b0),                                    // (terminated)
		.out_channel       ()                                         // (terminated)
	);

	Computer_System_DMA_1 dma_1 (
		.clk                  (system_pll_sys_clk_clk),                                      //                      clk.clk
		.reset                (rst_controller_reset_out_reset),                              //                    reset.reset
		.master_address       (dma_1_avalon_dma_master_address),                             //        avalon_dma_master.address
		.master_waitrequest   (dma_1_avalon_dma_master_waitrequest),                         //                         .waitrequest
		.master_arbiterlock   (dma_1_avalon_dma_master_lock),                                //                         .lock
		.master_read          (dma_1_avalon_dma_master_read),                                //                         .read
		.master_readdata      (dma_1_avalon_dma_master_readdata),                            //                         .readdata
		.master_readdatavalid (dma_1_avalon_dma_master_readdatavalid),                       //                         .readdatavalid
		.slave_address        (mm_interconnect_2_dma_1_avalon_dma_control_slave_address),    // avalon_dma_control_slave.address
		.slave_byteenable     (mm_interconnect_2_dma_1_avalon_dma_control_slave_byteenable), //                         .byteenable
		.slave_read           (mm_interconnect_2_dma_1_avalon_dma_control_slave_read),       //                         .read
		.slave_write          (mm_interconnect_2_dma_1_avalon_dma_control_slave_write),      //                         .write
		.slave_writedata      (mm_interconnect_2_dma_1_avalon_dma_control_slave_writedata),  //                         .writedata
		.slave_readdata       (mm_interconnect_2_dma_1_avalon_dma_control_slave_readdata),   //                         .readdata
		.stream_ready         (dma_1_avalon_pixel_source_ready),                             //      avalon_pixel_source.ready
		.stream_data          (dma_1_avalon_pixel_source_data),                              //                         .data
		.stream_startofpacket (dma_1_avalon_pixel_source_startofpacket),                     //                         .startofpacket
		.stream_endofpacket   (dma_1_avalon_pixel_source_endofpacket),                       //                         .endofpacket
		.stream_valid         (dma_1_avalon_pixel_source_valid)                              //                         .valid
	);

	Computer_System_DMA_1 dma_2 (
		.clk                  (system_pll_sys_clk_clk),                                      //                      clk.clk
		.reset                (rst_controller_reset_out_reset),                              //                    reset.reset
		.master_address       (dma_2_avalon_dma_master_address),                             //        avalon_dma_master.address
		.master_waitrequest   (dma_2_avalon_dma_master_waitrequest),                         //                         .waitrequest
		.master_arbiterlock   (dma_2_avalon_dma_master_lock),                                //                         .lock
		.master_read          (dma_2_avalon_dma_master_read),                                //                         .read
		.master_readdata      (dma_2_avalon_dma_master_readdata),                            //                         .readdata
		.master_readdatavalid (dma_2_avalon_dma_master_readdatavalid),                       //                         .readdatavalid
		.slave_address        (mm_interconnect_2_dma_2_avalon_dma_control_slave_address),    // avalon_dma_control_slave.address
		.slave_byteenable     (mm_interconnect_2_dma_2_avalon_dma_control_slave_byteenable), //                         .byteenable
		.slave_read           (mm_interconnect_2_dma_2_avalon_dma_control_slave_read),       //                         .read
		.slave_write          (mm_interconnect_2_dma_2_avalon_dma_control_slave_write),      //                         .write
		.slave_writedata      (mm_interconnect_2_dma_2_avalon_dma_control_slave_writedata),  //                         .writedata
		.slave_readdata       (mm_interconnect_2_dma_2_avalon_dma_control_slave_readdata),   //                         .readdata
		.stream_ready         (dma_2_avalon_pixel_source_ready),                             //      avalon_pixel_source.ready
		.stream_data          (dma_2_avalon_pixel_source_data),                              //                         .data
		.stream_startofpacket (dma_2_avalon_pixel_source_startofpacket),                     //                         .startofpacket
		.stream_endofpacket   (dma_2_avalon_pixel_source_endofpacket),                       //                         .endofpacket
		.stream_valid         (dma_2_avalon_pixel_source_valid)                              //                         .valid
	);

	Computer_System_DMA_WRITE dma_write (
		.clk                  (system_pll_sys_clk_clk),                                          //                      clk.clk
		.reset                (rst_controller_reset_out_reset),                                  //                    reset.reset
		.stream_data          (fusion_data_source_data),                                         //          avalon_dma_sink.data
		.stream_startofpacket (fusion_data_source_startofpacket),                                //                         .startofpacket
		.stream_endofpacket   (fusion_data_source_endofpacket),                                  //                         .endofpacket
		.stream_valid         (fusion_data_source_valid),                                        //                         .valid
		.stream_ready         (fusion_data_source_ready),                                        //                         .ready
		.slave_address        (mm_interconnect_2_dma_write_avalon_dma_control_slave_address),    // avalon_dma_control_slave.address
		.slave_byteenable     (mm_interconnect_2_dma_write_avalon_dma_control_slave_byteenable), //                         .byteenable
		.slave_read           (mm_interconnect_2_dma_write_avalon_dma_control_slave_read),       //                         .read
		.slave_write          (mm_interconnect_2_dma_write_avalon_dma_control_slave_write),      //                         .write
		.slave_writedata      (mm_interconnect_2_dma_write_avalon_dma_control_slave_writedata),  //                         .writedata
		.slave_readdata       (mm_interconnect_2_dma_write_avalon_dma_control_slave_readdata),   //                         .readdata
		.master_address       (dma_write_avalon_dma_master_address),                             //        avalon_dma_master.address
		.master_waitrequest   (dma_write_avalon_dma_master_waitrequest),                         //                         .waitrequest
		.master_write         (dma_write_avalon_dma_master_write),                               //                         .write
		.master_writedata     (dma_write_avalon_dma_master_writedata)                            //                         .writedata
	);

	localedgepreserve fusion (
		.reset        (rst_controller_reset_out_reset),                //       reset.reset
		.Clock        (system_pll_sys_clk_clk),                        //       clock.clk
		.sink1_data   (padding_1_avalon_clipper_source_data),          //  data1_sink.data
		.sink1_eop    (padding_1_avalon_clipper_source_endofpacket),   //            .endofpacket
		.sink1_ready  (padding_1_avalon_clipper_source_ready),         //            .ready
		.sink1_sop    (padding_1_avalon_clipper_source_startofpacket), //            .startofpacket
		.sink1_valid  (padding_1_avalon_clipper_source_valid),         //            .valid
		.sink2_data   (padding_2_avalon_clipper_source_data),          //  data2_sink.data
		.sink2_eop    (padding_2_avalon_clipper_source_endofpacket),   //            .endofpacket
		.sink2_ready  (padding_2_avalon_clipper_source_ready),         //            .ready
		.sink2_sop    (padding_2_avalon_clipper_source_startofpacket), //            .startofpacket
		.sink2_valid  (padding_2_avalon_clipper_source_valid),         //            .valid
		.source_data  (fusion_data_source_data),                       // data_source.data
		.source_eop   (fusion_data_source_endofpacket),                //            .endofpacket
		.source_ready (fusion_data_source_ready),                      //            .ready
		.source_sop   (fusion_data_source_startofpacket),              //            .startofpacket
		.source_valid (fusion_data_source_valid)                       //            .valid
	);

	Computer_System_PADDING_1 padding_1 (
		.clk                      (system_pll_sys_clk_clk),                        //                   clk.clk
		.reset                    (rst_controller_reset_out_reset),                //                 reset.reset
		.stream_in_data           (buffer_1_out_data),                             //   avalon_clipper_sink.data
		.stream_in_startofpacket  (buffer_1_out_startofpacket),                    //                      .startofpacket
		.stream_in_endofpacket    (buffer_1_out_endofpacket),                      //                      .endofpacket
		.stream_in_valid          (buffer_1_out_valid),                            //                      .valid
		.stream_in_ready          (buffer_1_out_ready),                            //                      .ready
		.stream_out_ready         (padding_1_avalon_clipper_source_ready),         // avalon_clipper_source.ready
		.stream_out_data          (padding_1_avalon_clipper_source_data),          //                      .data
		.stream_out_startofpacket (padding_1_avalon_clipper_source_startofpacket), //                      .startofpacket
		.stream_out_endofpacket   (padding_1_avalon_clipper_source_endofpacket),   //                      .endofpacket
		.stream_out_valid         (padding_1_avalon_clipper_source_valid)          //                      .valid
	);

	Computer_System_PADDING_1 padding_2 (
		.clk                      (system_pll_sys_clk_clk),                        //                   clk.clk
		.reset                    (rst_controller_reset_out_reset),                //                 reset.reset
		.stream_in_data           (buffer_2_out_data),                             //   avalon_clipper_sink.data
		.stream_in_startofpacket  (buffer_2_out_startofpacket),                    //                      .startofpacket
		.stream_in_endofpacket    (buffer_2_out_endofpacket),                      //                      .endofpacket
		.stream_in_valid          (buffer_2_out_valid),                            //                      .valid
		.stream_in_ready          (buffer_2_out_ready),                            //                      .ready
		.stream_out_ready         (padding_2_avalon_clipper_source_ready),         // avalon_clipper_source.ready
		.stream_out_data          (padding_2_avalon_clipper_source_data),          //                      .data
		.stream_out_startofpacket (padding_2_avalon_clipper_source_startofpacket), //                      .startofpacket
		.stream_out_endofpacket   (padding_2_avalon_clipper_source_endofpacket),   //                      .endofpacket
		.stream_out_valid         (padding_2_avalon_clipper_source_valid)          //                      .valid
	);

	Computer_System_RAM ram (
		.address     (mm_interconnect_1_ram_s1_address),    //     s1.address
		.clken       (mm_interconnect_1_ram_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_1_ram_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_1_ram_s1_write),      //       .write
		.readdata    (mm_interconnect_1_ram_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_1_ram_s1_writedata),  //       .writedata
		.address2    (mm_interconnect_4_ram_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_4_ram_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_4_ram_s2_clken),      //       .clken
		.write2      (mm_interconnect_4_ram_s2_write),      //       .write
		.readdata2   (mm_interconnect_4_ram_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_4_ram_s2_writedata),  //       .writedata
		.clk         (system_pll_sys_clk_clk),              //   clk1.clk
		.reset       (rst_controller_reset_out_reset),      // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),  //       .reset_req
		.freeze      (1'b0)                                 // (terminated)
	);

	Computer_System_SYSTEM_PLL system_pll (
		.ref_clk_clk        (system_pll_ref_clk_clk),        //      ref_clk.clk
		.ref_reset_reset    (system_pll_ref_reset_reset),    //    ref_reset.reset
		.sys_clk_clk        (system_pll_sys_clk_clk),        //      sys_clk.clk
		.sdram_clk_clk      (),                              //    sdram_clk.clk
		.reset_source_reset (system_pll_reset_source_reset)  // reset_source.reset
	);

	Computer_System_VGA_PLL vga_pll (
		.refclk   (system_pll_sys_clk_clk),             //  refclk.clk
		.rst      (rst_controller_001_reset_out_reset), //   reset.reset
		.outclk_0 (vga_clk_clk),                        // outclk0.clk
		.locked   ()                                    // (terminated)
	);

	Computer_System_VGA_SUBSYSTEM vga_subsystem (
		.pixel_dma_control_slave_address    (mm_interconnect_3_vga_subsystem_pixel_dma_control_slave_address),    // pixel_dma_control_slave.address
		.pixel_dma_control_slave_byteenable (mm_interconnect_3_vga_subsystem_pixel_dma_control_slave_byteenable), //                        .byteenable
		.pixel_dma_control_slave_read       (mm_interconnect_3_vga_subsystem_pixel_dma_control_slave_read),       //                        .read
		.pixel_dma_control_slave_write      (mm_interconnect_3_vga_subsystem_pixel_dma_control_slave_write),      //                        .write
		.pixel_dma_control_slave_writedata  (mm_interconnect_3_vga_subsystem_pixel_dma_control_slave_writedata),  //                        .writedata
		.pixel_dma_control_slave_readdata   (mm_interconnect_3_vga_subsystem_pixel_dma_control_slave_readdata),   //                        .readdata
		.pixel_dma_master_readdatavalid     (vga_subsystem_pixel_dma_master_readdatavalid),                       //        pixel_dma_master.readdatavalid
		.pixel_dma_master_waitrequest       (vga_subsystem_pixel_dma_master_waitrequest),                         //                        .waitrequest
		.pixel_dma_master_address           (vga_subsystem_pixel_dma_master_address),                             //                        .address
		.pixel_dma_master_lock              (vga_subsystem_pixel_dma_master_lock),                                //                        .lock
		.pixel_dma_master_read              (vga_subsystem_pixel_dma_master_read),                                //                        .read
		.pixel_dma_master_readdata          (vga_subsystem_pixel_dma_master_readdata),                            //                        .readdata
		.sys_clk_clk                        (system_pll_sys_clk_clk),                                             //                 sys_clk.clk
		.sys_reset_reset_n                  (~rst_controller_002_reset_out_reset),                                //               sys_reset.reset_n
		.vga_CLK                            (vga_CLK),                                                            //                     vga.CLK
		.vga_HS                             (vga_HS),                                                             //                        .HS
		.vga_VS                             (vga_VS),                                                             //                        .VS
		.vga_BLANK                          (vga_BLANK),                                                          //                        .BLANK
		.vga_SYNC                           (vga_SYNC),                                                           //                        .SYNC
		.vga_R                              (vga_R),                                                              //                        .R
		.vga_G                              (vga_G),                                                              //                        .G
		.vga_B                              (vga_B),                                                              //                        .B
		.vga_pll_ref_clk_clk                (vga_pll_ref_clk_clk),                                                //         vga_pll_ref_clk.clk
		.vga_pll_ref_reset_reset            (vga_pll_ref_reset_reset)                                             //       vga_pll_ref_reset.reset
	);

	altera_up_avalon_video_dma_ctrl_addr_trans #(
		.ADDRESS_TRANSLATION_MASK (32'b11000000000000000000000000000000)
	) video_dma_address_translator (
		.clk                (system_pll_sys_clk_clk),                                           //  clock.clk
		.reset              (rst_controller_reset_out_reset),                                   //  reset.reset
		.slave_address      (mm_interconnect_2_video_dma_address_translator_slave_address),     //  slave.address
		.slave_byteenable   (mm_interconnect_2_video_dma_address_translator_slave_byteenable),  //       .byteenable
		.slave_read         (mm_interconnect_2_video_dma_address_translator_slave_read),        //       .read
		.slave_write        (mm_interconnect_2_video_dma_address_translator_slave_write),       //       .write
		.slave_writedata    (mm_interconnect_2_video_dma_address_translator_slave_writedata),   //       .writedata
		.slave_readdata     (mm_interconnect_2_video_dma_address_translator_slave_readdata),    //       .readdata
		.slave_waitrequest  (mm_interconnect_2_video_dma_address_translator_slave_waitrequest), //       .waitrequest
		.master_readdata    (video_dma_address_translator_master_readdata),                     // master.readdata
		.master_waitrequest (video_dma_address_translator_master_waitrequest),                  //       .waitrequest
		.master_address     (video_dma_address_translator_master_address),                      //       .address
		.master_byteenable  (video_dma_address_translator_master_byteenable),                   //       .byteenable
		.master_read        (video_dma_address_translator_master_read),                         //       .read
		.master_write       (video_dma_address_translator_master_write),                        //       .write
		.master_writedata   (video_dma_address_translator_master_writedata)                     //       .writedata
	);

	Computer_System_mm_interconnect_0 mm_interconnect_0 (
		.ARM_A9_HPS_f2h_axi_slave_awid                                         (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awid),    //                                        ARM_A9_HPS_f2h_axi_slave.awid
		.ARM_A9_HPS_f2h_axi_slave_awaddr                                       (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awaddr),  //                                                                .awaddr
		.ARM_A9_HPS_f2h_axi_slave_awlen                                        (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awlen),   //                                                                .awlen
		.ARM_A9_HPS_f2h_axi_slave_awsize                                       (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awsize),  //                                                                .awsize
		.ARM_A9_HPS_f2h_axi_slave_awburst                                      (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awburst), //                                                                .awburst
		.ARM_A9_HPS_f2h_axi_slave_awlock                                       (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awlock),  //                                                                .awlock
		.ARM_A9_HPS_f2h_axi_slave_awcache                                      (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awcache), //                                                                .awcache
		.ARM_A9_HPS_f2h_axi_slave_awprot                                       (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awprot),  //                                                                .awprot
		.ARM_A9_HPS_f2h_axi_slave_awuser                                       (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awuser),  //                                                                .awuser
		.ARM_A9_HPS_f2h_axi_slave_awvalid                                      (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awvalid), //                                                                .awvalid
		.ARM_A9_HPS_f2h_axi_slave_awready                                      (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awready), //                                                                .awready
		.ARM_A9_HPS_f2h_axi_slave_wid                                          (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_wid),     //                                                                .wid
		.ARM_A9_HPS_f2h_axi_slave_wdata                                        (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_wdata),   //                                                                .wdata
		.ARM_A9_HPS_f2h_axi_slave_wstrb                                        (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_wstrb),   //                                                                .wstrb
		.ARM_A9_HPS_f2h_axi_slave_wlast                                        (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_wlast),   //                                                                .wlast
		.ARM_A9_HPS_f2h_axi_slave_wvalid                                       (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_wvalid),  //                                                                .wvalid
		.ARM_A9_HPS_f2h_axi_slave_wready                                       (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_wready),  //                                                                .wready
		.ARM_A9_HPS_f2h_axi_slave_bid                                          (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_bid),     //                                                                .bid
		.ARM_A9_HPS_f2h_axi_slave_bresp                                        (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_bresp),   //                                                                .bresp
		.ARM_A9_HPS_f2h_axi_slave_bvalid                                       (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_bvalid),  //                                                                .bvalid
		.ARM_A9_HPS_f2h_axi_slave_bready                                       (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_bready),  //                                                                .bready
		.ARM_A9_HPS_f2h_axi_slave_arid                                         (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arid),    //                                                                .arid
		.ARM_A9_HPS_f2h_axi_slave_araddr                                       (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_araddr),  //                                                                .araddr
		.ARM_A9_HPS_f2h_axi_slave_arlen                                        (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arlen),   //                                                                .arlen
		.ARM_A9_HPS_f2h_axi_slave_arsize                                       (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arsize),  //                                                                .arsize
		.ARM_A9_HPS_f2h_axi_slave_arburst                                      (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arburst), //                                                                .arburst
		.ARM_A9_HPS_f2h_axi_slave_arlock                                       (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arlock),  //                                                                .arlock
		.ARM_A9_HPS_f2h_axi_slave_arcache                                      (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arcache), //                                                                .arcache
		.ARM_A9_HPS_f2h_axi_slave_arprot                                       (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arprot),  //                                                                .arprot
		.ARM_A9_HPS_f2h_axi_slave_aruser                                       (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_aruser),  //                                                                .aruser
		.ARM_A9_HPS_f2h_axi_slave_arvalid                                      (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arvalid), //                                                                .arvalid
		.ARM_A9_HPS_f2h_axi_slave_arready                                      (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arready), //                                                                .arready
		.ARM_A9_HPS_f2h_axi_slave_rid                                          (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_rid),     //                                                                .rid
		.ARM_A9_HPS_f2h_axi_slave_rdata                                        (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_rdata),   //                                                                .rdata
		.ARM_A9_HPS_f2h_axi_slave_rresp                                        (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_rresp),   //                                                                .rresp
		.ARM_A9_HPS_f2h_axi_slave_rlast                                        (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_rlast),   //                                                                .rlast
		.ARM_A9_HPS_f2h_axi_slave_rvalid                                       (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_rvalid),  //                                                                .rvalid
		.ARM_A9_HPS_f2h_axi_slave_rready                                       (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_rready),  //                                                                .rready
		.SYSTEM_PLL_sys_clk_clk                                                (system_pll_sys_clk_clk),                             //                                              SYSTEM_PLL_sys_clk.clk
		.ARM_A9_HPS_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset_reset (rst_controller_003_reset_out_reset),                 // ARM_A9_HPS_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset.reset
		.DMA_1_reset_reset_bridge_in_reset_reset                               (rst_controller_reset_out_reset),                     //                               DMA_1_reset_reset_bridge_in_reset.reset
		.DMA_1_avalon_dma_master_address                                       (dma_1_avalon_dma_master_address),                    //                                         DMA_1_avalon_dma_master.address
		.DMA_1_avalon_dma_master_waitrequest                                   (dma_1_avalon_dma_master_waitrequest),                //                                                                .waitrequest
		.DMA_1_avalon_dma_master_read                                          (dma_1_avalon_dma_master_read),                       //                                                                .read
		.DMA_1_avalon_dma_master_readdata                                      (dma_1_avalon_dma_master_readdata),                   //                                                                .readdata
		.DMA_1_avalon_dma_master_readdatavalid                                 (dma_1_avalon_dma_master_readdatavalid),              //                                                                .readdatavalid
		.DMA_1_avalon_dma_master_lock                                          (dma_1_avalon_dma_master_lock),                       //                                                                .lock
		.DMA_2_avalon_dma_master_address                                       (dma_2_avalon_dma_master_address),                    //                                         DMA_2_avalon_dma_master.address
		.DMA_2_avalon_dma_master_waitrequest                                   (dma_2_avalon_dma_master_waitrequest),                //                                                                .waitrequest
		.DMA_2_avalon_dma_master_read                                          (dma_2_avalon_dma_master_read),                       //                                                                .read
		.DMA_2_avalon_dma_master_readdata                                      (dma_2_avalon_dma_master_readdata),                   //                                                                .readdata
		.DMA_2_avalon_dma_master_readdatavalid                                 (dma_2_avalon_dma_master_readdatavalid),              //                                                                .readdatavalid
		.DMA_2_avalon_dma_master_lock                                          (dma_2_avalon_dma_master_lock)                        //                                                                .lock
	);

	Computer_System_mm_interconnect_1 mm_interconnect_1 (
		.SYSTEM_PLL_sys_clk_clk                      (system_pll_sys_clk_clk),                  //                    SYSTEM_PLL_sys_clk.clk
		.DMA_WRITE_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),          // DMA_WRITE_reset_reset_bridge_in_reset.reset
		.DMA_WRITE_avalon_dma_master_address         (dma_write_avalon_dma_master_address),     //           DMA_WRITE_avalon_dma_master.address
		.DMA_WRITE_avalon_dma_master_waitrequest     (dma_write_avalon_dma_master_waitrequest), //                                      .waitrequest
		.DMA_WRITE_avalon_dma_master_write           (dma_write_avalon_dma_master_write),       //                                      .write
		.DMA_WRITE_avalon_dma_master_writedata       (dma_write_avalon_dma_master_writedata),   //                                      .writedata
		.RAM_s1_address                              (mm_interconnect_1_ram_s1_address),        //                                RAM_s1.address
		.RAM_s1_write                                (mm_interconnect_1_ram_s1_write),          //                                      .write
		.RAM_s1_readdata                             (mm_interconnect_1_ram_s1_readdata),       //                                      .readdata
		.RAM_s1_writedata                            (mm_interconnect_1_ram_s1_writedata),      //                                      .writedata
		.RAM_s1_chipselect                           (mm_interconnect_1_ram_s1_chipselect),     //                                      .chipselect
		.RAM_s1_clken                                (mm_interconnect_1_ram_s1_clken)           //                                      .clken
	);

	Computer_System_mm_interconnect_2 mm_interconnect_2 (
		.ARM_A9_HPS_h2f_lw_axi_master_awid                                        (arm_a9_hps_h2f_lw_axi_master_awid),                                //                                       ARM_A9_HPS_h2f_lw_axi_master.awid
		.ARM_A9_HPS_h2f_lw_axi_master_awaddr                                      (arm_a9_hps_h2f_lw_axi_master_awaddr),                              //                                                                   .awaddr
		.ARM_A9_HPS_h2f_lw_axi_master_awlen                                       (arm_a9_hps_h2f_lw_axi_master_awlen),                               //                                                                   .awlen
		.ARM_A9_HPS_h2f_lw_axi_master_awsize                                      (arm_a9_hps_h2f_lw_axi_master_awsize),                              //                                                                   .awsize
		.ARM_A9_HPS_h2f_lw_axi_master_awburst                                     (arm_a9_hps_h2f_lw_axi_master_awburst),                             //                                                                   .awburst
		.ARM_A9_HPS_h2f_lw_axi_master_awlock                                      (arm_a9_hps_h2f_lw_axi_master_awlock),                              //                                                                   .awlock
		.ARM_A9_HPS_h2f_lw_axi_master_awcache                                     (arm_a9_hps_h2f_lw_axi_master_awcache),                             //                                                                   .awcache
		.ARM_A9_HPS_h2f_lw_axi_master_awprot                                      (arm_a9_hps_h2f_lw_axi_master_awprot),                              //                                                                   .awprot
		.ARM_A9_HPS_h2f_lw_axi_master_awvalid                                     (arm_a9_hps_h2f_lw_axi_master_awvalid),                             //                                                                   .awvalid
		.ARM_A9_HPS_h2f_lw_axi_master_awready                                     (arm_a9_hps_h2f_lw_axi_master_awready),                             //                                                                   .awready
		.ARM_A9_HPS_h2f_lw_axi_master_wid                                         (arm_a9_hps_h2f_lw_axi_master_wid),                                 //                                                                   .wid
		.ARM_A9_HPS_h2f_lw_axi_master_wdata                                       (arm_a9_hps_h2f_lw_axi_master_wdata),                               //                                                                   .wdata
		.ARM_A9_HPS_h2f_lw_axi_master_wstrb                                       (arm_a9_hps_h2f_lw_axi_master_wstrb),                               //                                                                   .wstrb
		.ARM_A9_HPS_h2f_lw_axi_master_wlast                                       (arm_a9_hps_h2f_lw_axi_master_wlast),                               //                                                                   .wlast
		.ARM_A9_HPS_h2f_lw_axi_master_wvalid                                      (arm_a9_hps_h2f_lw_axi_master_wvalid),                              //                                                                   .wvalid
		.ARM_A9_HPS_h2f_lw_axi_master_wready                                      (arm_a9_hps_h2f_lw_axi_master_wready),                              //                                                                   .wready
		.ARM_A9_HPS_h2f_lw_axi_master_bid                                         (arm_a9_hps_h2f_lw_axi_master_bid),                                 //                                                                   .bid
		.ARM_A9_HPS_h2f_lw_axi_master_bresp                                       (arm_a9_hps_h2f_lw_axi_master_bresp),                               //                                                                   .bresp
		.ARM_A9_HPS_h2f_lw_axi_master_bvalid                                      (arm_a9_hps_h2f_lw_axi_master_bvalid),                              //                                                                   .bvalid
		.ARM_A9_HPS_h2f_lw_axi_master_bready                                      (arm_a9_hps_h2f_lw_axi_master_bready),                              //                                                                   .bready
		.ARM_A9_HPS_h2f_lw_axi_master_arid                                        (arm_a9_hps_h2f_lw_axi_master_arid),                                //                                                                   .arid
		.ARM_A9_HPS_h2f_lw_axi_master_araddr                                      (arm_a9_hps_h2f_lw_axi_master_araddr),                              //                                                                   .araddr
		.ARM_A9_HPS_h2f_lw_axi_master_arlen                                       (arm_a9_hps_h2f_lw_axi_master_arlen),                               //                                                                   .arlen
		.ARM_A9_HPS_h2f_lw_axi_master_arsize                                      (arm_a9_hps_h2f_lw_axi_master_arsize),                              //                                                                   .arsize
		.ARM_A9_HPS_h2f_lw_axi_master_arburst                                     (arm_a9_hps_h2f_lw_axi_master_arburst),                             //                                                                   .arburst
		.ARM_A9_HPS_h2f_lw_axi_master_arlock                                      (arm_a9_hps_h2f_lw_axi_master_arlock),                              //                                                                   .arlock
		.ARM_A9_HPS_h2f_lw_axi_master_arcache                                     (arm_a9_hps_h2f_lw_axi_master_arcache),                             //                                                                   .arcache
		.ARM_A9_HPS_h2f_lw_axi_master_arprot                                      (arm_a9_hps_h2f_lw_axi_master_arprot),                              //                                                                   .arprot
		.ARM_A9_HPS_h2f_lw_axi_master_arvalid                                     (arm_a9_hps_h2f_lw_axi_master_arvalid),                             //                                                                   .arvalid
		.ARM_A9_HPS_h2f_lw_axi_master_arready                                     (arm_a9_hps_h2f_lw_axi_master_arready),                             //                                                                   .arready
		.ARM_A9_HPS_h2f_lw_axi_master_rid                                         (arm_a9_hps_h2f_lw_axi_master_rid),                                 //                                                                   .rid
		.ARM_A9_HPS_h2f_lw_axi_master_rdata                                       (arm_a9_hps_h2f_lw_axi_master_rdata),                               //                                                                   .rdata
		.ARM_A9_HPS_h2f_lw_axi_master_rresp                                       (arm_a9_hps_h2f_lw_axi_master_rresp),                               //                                                                   .rresp
		.ARM_A9_HPS_h2f_lw_axi_master_rlast                                       (arm_a9_hps_h2f_lw_axi_master_rlast),                               //                                                                   .rlast
		.ARM_A9_HPS_h2f_lw_axi_master_rvalid                                      (arm_a9_hps_h2f_lw_axi_master_rvalid),                              //                                                                   .rvalid
		.ARM_A9_HPS_h2f_lw_axi_master_rready                                      (arm_a9_hps_h2f_lw_axi_master_rready),                              //                                                                   .rready
		.SYSTEM_PLL_sys_clk_clk                                                   (system_pll_sys_clk_clk),                                           //                                                 SYSTEM_PLL_sys_clk.clk
		.ARM_A9_HPS_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_003_reset_out_reset),                               // ARM_A9_HPS_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.DMA_1_reset_reset_bridge_in_reset_reset                                  (rst_controller_reset_out_reset),                                   //                                  DMA_1_reset_reset_bridge_in_reset.reset
		.DMA_1_avalon_dma_control_slave_address                                   (mm_interconnect_2_dma_1_avalon_dma_control_slave_address),         //                                     DMA_1_avalon_dma_control_slave.address
		.DMA_1_avalon_dma_control_slave_write                                     (mm_interconnect_2_dma_1_avalon_dma_control_slave_write),           //                                                                   .write
		.DMA_1_avalon_dma_control_slave_read                                      (mm_interconnect_2_dma_1_avalon_dma_control_slave_read),            //                                                                   .read
		.DMA_1_avalon_dma_control_slave_readdata                                  (mm_interconnect_2_dma_1_avalon_dma_control_slave_readdata),        //                                                                   .readdata
		.DMA_1_avalon_dma_control_slave_writedata                                 (mm_interconnect_2_dma_1_avalon_dma_control_slave_writedata),       //                                                                   .writedata
		.DMA_1_avalon_dma_control_slave_byteenable                                (mm_interconnect_2_dma_1_avalon_dma_control_slave_byteenable),      //                                                                   .byteenable
		.DMA_2_avalon_dma_control_slave_address                                   (mm_interconnect_2_dma_2_avalon_dma_control_slave_address),         //                                     DMA_2_avalon_dma_control_slave.address
		.DMA_2_avalon_dma_control_slave_write                                     (mm_interconnect_2_dma_2_avalon_dma_control_slave_write),           //                                                                   .write
		.DMA_2_avalon_dma_control_slave_read                                      (mm_interconnect_2_dma_2_avalon_dma_control_slave_read),            //                                                                   .read
		.DMA_2_avalon_dma_control_slave_readdata                                  (mm_interconnect_2_dma_2_avalon_dma_control_slave_readdata),        //                                                                   .readdata
		.DMA_2_avalon_dma_control_slave_writedata                                 (mm_interconnect_2_dma_2_avalon_dma_control_slave_writedata),       //                                                                   .writedata
		.DMA_2_avalon_dma_control_slave_byteenable                                (mm_interconnect_2_dma_2_avalon_dma_control_slave_byteenable),      //                                                                   .byteenable
		.DMA_WRITE_avalon_dma_control_slave_address                               (mm_interconnect_2_dma_write_avalon_dma_control_slave_address),     //                                 DMA_WRITE_avalon_dma_control_slave.address
		.DMA_WRITE_avalon_dma_control_slave_write                                 (mm_interconnect_2_dma_write_avalon_dma_control_slave_write),       //                                                                   .write
		.DMA_WRITE_avalon_dma_control_slave_read                                  (mm_interconnect_2_dma_write_avalon_dma_control_slave_read),        //                                                                   .read
		.DMA_WRITE_avalon_dma_control_slave_readdata                              (mm_interconnect_2_dma_write_avalon_dma_control_slave_readdata),    //                                                                   .readdata
		.DMA_WRITE_avalon_dma_control_slave_writedata                             (mm_interconnect_2_dma_write_avalon_dma_control_slave_writedata),   //                                                                   .writedata
		.DMA_WRITE_avalon_dma_control_slave_byteenable                            (mm_interconnect_2_dma_write_avalon_dma_control_slave_byteenable),  //                                                                   .byteenable
		.VIDEO_DMA_ADDRESS_TRANSLATOR_slave_address                               (mm_interconnect_2_video_dma_address_translator_slave_address),     //                                 VIDEO_DMA_ADDRESS_TRANSLATOR_slave.address
		.VIDEO_DMA_ADDRESS_TRANSLATOR_slave_write                                 (mm_interconnect_2_video_dma_address_translator_slave_write),       //                                                                   .write
		.VIDEO_DMA_ADDRESS_TRANSLATOR_slave_read                                  (mm_interconnect_2_video_dma_address_translator_slave_read),        //                                                                   .read
		.VIDEO_DMA_ADDRESS_TRANSLATOR_slave_readdata                              (mm_interconnect_2_video_dma_address_translator_slave_readdata),    //                                                                   .readdata
		.VIDEO_DMA_ADDRESS_TRANSLATOR_slave_writedata                             (mm_interconnect_2_video_dma_address_translator_slave_writedata),   //                                                                   .writedata
		.VIDEO_DMA_ADDRESS_TRANSLATOR_slave_byteenable                            (mm_interconnect_2_video_dma_address_translator_slave_byteenable),  //                                                                   .byteenable
		.VIDEO_DMA_ADDRESS_TRANSLATOR_slave_waitrequest                           (mm_interconnect_2_video_dma_address_translator_slave_waitrequest)  //                                                                   .waitrequest
	);

	Computer_System_mm_interconnect_3 mm_interconnect_3 (
		.SYSTEM_PLL_sys_clk_clk                                         (system_pll_sys_clk_clk),                                             //                                       SYSTEM_PLL_sys_clk.clk
		.VGA_SUBSYSTEM_sys_reset_reset_bridge_in_reset_reset            (rst_controller_reset_out_reset),                                     //            VGA_SUBSYSTEM_sys_reset_reset_bridge_in_reset.reset
		.VIDEO_DMA_ADDRESS_TRANSLATOR_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                                     // VIDEO_DMA_ADDRESS_TRANSLATOR_reset_reset_bridge_in_reset.reset
		.VIDEO_DMA_ADDRESS_TRANSLATOR_master_address                    (video_dma_address_translator_master_address),                        //                      VIDEO_DMA_ADDRESS_TRANSLATOR_master.address
		.VIDEO_DMA_ADDRESS_TRANSLATOR_master_waitrequest                (video_dma_address_translator_master_waitrequest),                    //                                                         .waitrequest
		.VIDEO_DMA_ADDRESS_TRANSLATOR_master_byteenable                 (video_dma_address_translator_master_byteenable),                     //                                                         .byteenable
		.VIDEO_DMA_ADDRESS_TRANSLATOR_master_read                       (video_dma_address_translator_master_read),                           //                                                         .read
		.VIDEO_DMA_ADDRESS_TRANSLATOR_master_readdata                   (video_dma_address_translator_master_readdata),                       //                                                         .readdata
		.VIDEO_DMA_ADDRESS_TRANSLATOR_master_write                      (video_dma_address_translator_master_write),                          //                                                         .write
		.VIDEO_DMA_ADDRESS_TRANSLATOR_master_writedata                  (video_dma_address_translator_master_writedata),                      //                                                         .writedata
		.VGA_SUBSYSTEM_pixel_dma_control_slave_address                  (mm_interconnect_3_vga_subsystem_pixel_dma_control_slave_address),    //                    VGA_SUBSYSTEM_pixel_dma_control_slave.address
		.VGA_SUBSYSTEM_pixel_dma_control_slave_write                    (mm_interconnect_3_vga_subsystem_pixel_dma_control_slave_write),      //                                                         .write
		.VGA_SUBSYSTEM_pixel_dma_control_slave_read                     (mm_interconnect_3_vga_subsystem_pixel_dma_control_slave_read),       //                                                         .read
		.VGA_SUBSYSTEM_pixel_dma_control_slave_readdata                 (mm_interconnect_3_vga_subsystem_pixel_dma_control_slave_readdata),   //                                                         .readdata
		.VGA_SUBSYSTEM_pixel_dma_control_slave_writedata                (mm_interconnect_3_vga_subsystem_pixel_dma_control_slave_writedata),  //                                                         .writedata
		.VGA_SUBSYSTEM_pixel_dma_control_slave_byteenable               (mm_interconnect_3_vga_subsystem_pixel_dma_control_slave_byteenable)  //                                                         .byteenable
	);

	Computer_System_mm_interconnect_4 mm_interconnect_4 (
		.SYSTEM_PLL_sys_clk_clk                              (system_pll_sys_clk_clk),                       //                            SYSTEM_PLL_sys_clk.clk
		.RAM_reset1_reset_bridge_in_reset_reset              (rst_controller_reset_out_reset),               //              RAM_reset1_reset_bridge_in_reset.reset
		.VGA_SUBSYSTEM_sys_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),               // VGA_SUBSYSTEM_sys_reset_reset_bridge_in_reset.reset
		.VGA_SUBSYSTEM_pixel_dma_master_address              (vga_subsystem_pixel_dma_master_address),       //                VGA_SUBSYSTEM_pixel_dma_master.address
		.VGA_SUBSYSTEM_pixel_dma_master_waitrequest          (vga_subsystem_pixel_dma_master_waitrequest),   //                                              .waitrequest
		.VGA_SUBSYSTEM_pixel_dma_master_read                 (vga_subsystem_pixel_dma_master_read),          //                                              .read
		.VGA_SUBSYSTEM_pixel_dma_master_readdata             (vga_subsystem_pixel_dma_master_readdata),      //                                              .readdata
		.VGA_SUBSYSTEM_pixel_dma_master_readdatavalid        (vga_subsystem_pixel_dma_master_readdatavalid), //                                              .readdatavalid
		.VGA_SUBSYSTEM_pixel_dma_master_lock                 (vga_subsystem_pixel_dma_master_lock),          //                                              .lock
		.RAM_s2_address                                      (mm_interconnect_4_ram_s2_address),             //                                        RAM_s2.address
		.RAM_s2_write                                        (mm_interconnect_4_ram_s2_write),               //                                              .write
		.RAM_s2_readdata                                     (mm_interconnect_4_ram_s2_readdata),            //                                              .readdata
		.RAM_s2_writedata                                    (mm_interconnect_4_ram_s2_writedata),           //                                              .writedata
		.RAM_s2_chipselect                                   (mm_interconnect_4_ram_s2_chipselect),          //                                              .chipselect
		.RAM_s2_clken                                        (mm_interconnect_4_ram_s2_clken)                //                                              .clken
	);

	Computer_System_irq_mapper irq_mapper (
		.clk        (),                        //       clk.clk
		.reset      (),                        // clk_reset.reset
		.sender_irq (arm_a9_hps_f2h_irq0_irq)  //    sender.irq
	);

	Computer_System_irq_mapper irq_mapper_001 (
		.clk        (),                        //       clk.clk
		.reset      (),                        // clk_reset.reset
		.sender_irq (arm_a9_hps_f2h_irq1_irq)  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~arm_a9_hps_h2f_reset_reset),        // reset_in0.reset
		.reset_in1      (system_pll_reset_source_reset),      // reset_in1.reset
		.clk            (system_pll_sys_clk_clk),             //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~arm_a9_hps_h2f_reset_reset),        // reset_in0.reset
		.reset_in1      (system_pll_reset_source_reset),      // reset_in1.reset
		.clk            (),                                   //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~arm_a9_hps_h2f_reset_reset),        // reset_in0.reset
		.reset_in1      (system_pll_reset_source_reset),      // reset_in1.reset
		.clk            (),                                   //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~arm_a9_hps_h2f_reset_reset),        // reset_in0.reset
		.clk            (system_pll_sys_clk_clk),             //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
