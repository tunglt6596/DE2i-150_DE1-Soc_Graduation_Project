-- gaussian_ip_GN_gaussian_ip_Fusion.vhd

-- Generated using ACDS version 17.1 590

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity gaussian_ip_GN_gaussian_ip_Fusion is
	port (
		sof_out   : out std_logic_vector(0 downto 0);                    --   sof_out.wire
		pixel2_in : in  std_logic_vector(7 downto 0) := (others => '0'); -- pixel2_in.wire
		sof1_in   : in  std_logic                    := '0';             --   sof1_in.wire
		ready2_in : out std_logic;                                       -- ready2_in.wire
		valid1_in : in  std_logic                    := '0';             -- valid1_in.wire
		valid_out : out std_logic_vector(0 downto 0);                    -- valid_out.wire
		eof1_in   : in  std_logic                    := '0';             --   eof1_in.wire
		pixel1_in : in  std_logic_vector(7 downto 0) := (others => '0'); -- pixel1_in.wire
		eof_out   : out std_logic_vector(0 downto 0);                    --   eof_out.wire
		Clock     : in  std_logic                    := '0';             --     Clock.clk
		reset     : in  std_logic                    := '0';             --          .reset
		pixel_out : out std_logic_vector(9 downto 0)                     -- pixel_out.wire
	);
end entity gaussian_ip_GN_gaussian_ip_Fusion;

architecture rtl of gaussian_ip_GN_gaussian_ip_Fusion is
	component alt_dspbuilder_clock_GNQFU4PUDH is
		port (
			aclr      : in  std_logic := 'X'; -- reset
			aclr_n    : in  std_logic := 'X'; -- reset_n
			aclr_out  : out std_logic;        -- reset
			clock     : in  std_logic := 'X'; -- clk
			clock_out : out std_logic         -- clk
		);
	end component alt_dspbuilder_clock_GNQFU4PUDH;

	component alt_dspbuilder_port_GNXAOKDYKC is
		port (
			input  : in  std_logic_vector(0 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(0 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNXAOKDYKC;

	component alt_dspbuilder_port_GNA5S4SQDN is
		port (
			input  : in  std_logic_vector(7 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(7 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNA5S4SQDN;

	component alt_dspbuilder_multiplexer_GNWZZP2IFI is
		generic (
			number_inputs          : natural  := 4;
			pipeline               : natural  := 0;
			width                  : positive := 8;
			HDLTYPE                : string   := "STD_LOGIC_VECTOR";
			use_one_hot_select_bus : natural  := 0
		);
		port (
			clock     : in  std_logic                    := 'X';             -- clk
			aclr      : in  std_logic                    := 'X';             -- reset
			sel       : in  std_logic_vector(0 downto 0) := (others => 'X'); -- wire
			result    : out std_logic_vector(9 downto 0);                    -- wire
			ena       : in  std_logic                    := 'X';             -- wire
			user_aclr : in  std_logic                    := 'X';             -- wire
			in0       : in  std_logic_vector(9 downto 0) := (others => 'X'); -- wire
			in1       : in  std_logic_vector(9 downto 0) := (others => 'X')  -- wire
		);
	end component alt_dspbuilder_multiplexer_GNWZZP2IFI;

	component alt_dspbuilder_gnd_GN is
		port (
			output : out std_logic   -- wire
		);
	end component alt_dspbuilder_gnd_GN;

	component alt_dspbuilder_vcc_GN is
		port (
			output : out std_logic   -- wire
		);
	end component alt_dspbuilder_vcc_GN;

	component alt_dspbuilder_port_GN37ALZBS4 is
		port (
			input  : in  std_logic := 'X'; -- wire
			output : out std_logic         -- wire
		);
	end component alt_dspbuilder_port_GN37ALZBS4;

	component alt_dspbuilder_constant_GN6SFEINY6 is
		generic (
			BitPattern : string  := "0000";
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(1 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GN6SFEINY6;

	component alt_dspbuilder_pipelined_adder_GN4HTUTWRG is
		generic (
			pipeline : integer := 0;
			width    : natural := 0
		);
		port (
			aclr      : in  std_logic                          := 'X';             -- clk
			add_sub   : in  std_logic                          := 'X';             -- wire
			cin       : in  std_logic                          := 'X';             -- wire
			clock     : in  std_logic                          := 'X';             -- clk
			cout      : out std_logic;                                             -- wire
			dataa     : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			datab     : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			ena       : in  std_logic                          := 'X';             -- wire
			result    : out std_logic_vector(width-1 downto 0);                    -- wire
			user_aclr : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_pipelined_adder_GN4HTUTWRG;

	component alt_dspbuilder_comparator_GN is
		generic (
			Operator  : string  := "Altaeb";
			lpm_width : natural := 8
		);
		port (
			clock  : in  std_logic                              := 'X';             -- clk
			dataa  : in  std_logic_vector(lpm_width-1 downto 0) := (others => 'X'); -- wire
			datab  : in  std_logic_vector(lpm_width-1 downto 0) := (others => 'X'); -- wire
			result : out std_logic;                                                 -- wire
			sclr   : in  std_logic                              := 'X'              -- clk
		);
	end component alt_dspbuilder_comparator_GN;

	component alt_dspbuilder_memdelay_GNR55NYJWV is
		generic (
			RAMTYPE : string   := "AUTO";
			WIDTH   : positive := 8;
			DELAY   : positive := 1
		);
		port (
			aclr      : in  std_logic                          := 'X';             -- clk
			clock     : in  std_logic                          := 'X';             -- clk
			ena       : in  std_logic                          := 'X';             -- wire
			input     : in  std_logic_vector(WIDTH-1 downto 0) := (others => 'X'); -- wire
			output    : out std_logic_vector(WIDTH-1 downto 0);                    -- wire
			user_aclr : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_memdelay_GNR55NYJWV;

	component alt_dspbuilder_constant_GNC5NOVIJT is
		generic (
			BitPattern : string  := "0000";
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(7 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GNC5NOVIJT;

	component alt_dspbuilder_constant_GNSVSRQZMI is
		generic (
			BitPattern : string  := "0000";
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(7 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GNSVSRQZMI;

	component alt_dspbuilder_constant_GN5IRMZXKK is
		generic (
			BitPattern : string  := "0000";
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(9 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GN5IRMZXKK;

	component alt_dspbuilder_bus_concat_GNKLOJ6ING is
		generic (
			widthA : natural := 8;
			widthB : natural := 8
		);
		port (
			a      : in  std_logic_vector(widthA-1 downto 0)        := (others => 'X'); -- wire
			aclr   : in  std_logic                                  := 'X';             -- clk
			b      : in  std_logic_vector(widthB-1 downto 0)        := (others => 'X'); -- wire
			clock  : in  std_logic                                  := 'X';             -- clk
			output : out std_logic_vector(widthA+widthB-1 downto 0)                     -- wire
		);
	end component alt_dspbuilder_bus_concat_GNKLOJ6ING;

	component alt_dspbuilder_constant_GNK57PM5EK is
		generic (
			BitPattern : string  := "0000";
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(9 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GNK57PM5EK;

	component alt_dspbuilder_memdelay_GNT3M75IMA is
		generic (
			RAMTYPE : string   := "AUTO";
			WIDTH   : positive := 8;
			DELAY   : positive := 1
		);
		port (
			aclr      : in  std_logic                          := 'X';             -- clk
			clock     : in  std_logic                          := 'X';             -- clk
			ena       : in  std_logic                          := 'X';             -- wire
			input     : in  std_logic_vector(WIDTH-1 downto 0) := (others => 'X'); -- wire
			output    : out std_logic_vector(WIDTH-1 downto 0);                    -- wire
			user_aclr : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_memdelay_GNT3M75IMA;

	component alt_dspbuilder_port_GNSSYS4J5R is
		port (
			input  : in  std_logic_vector(9 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(9 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNSSYS4J5R;

	component gaussian_ip_GN_gaussian_ip_Fusion_Decomposition_3 is
		port (
			sof_in    : in  std_logic                    := 'X';             -- wire
			sof_out   : out std_logic;                                       -- wire
			Clock     : in  std_logic                    := 'X';             -- clk
			reset     : in  std_logic                    := 'X';             -- reset
			eof_in    : in  std_logic                    := 'X';             -- wire
			eof_out   : out std_logic;                                       -- wire
			valid_in  : in  std_logic                    := 'X';             -- wire
			diff_out  : out std_logic_vector(9 downto 0);                    -- wire
			valid_out : out std_logic;                                       -- wire
			diff_in   : in  std_logic_vector(9 downto 0) := (others => 'X'); -- wire
			pixel_out : out std_logic_vector(7 downto 0);                    -- wire
			pixel_in  : in  std_logic_vector(7 downto 0) := (others => 'X')  -- wire
		);
	end component gaussian_ip_GN_gaussian_ip_Fusion_Decomposition_3;

	component gaussian_ip_GN_gaussian_ip_Fusion_Decomposition_1 is
		port (
			valid_in  : in  std_logic                    := 'X';             -- wire
			valid_out : out std_logic;                                       -- wire
			pixel_out : out std_logic_vector(7 downto 0);                    -- wire
			diff_out  : out std_logic_vector(9 downto 0);                    -- wire
			eof_out   : out std_logic;                                       -- wire
			sof_in    : in  std_logic                    := 'X';             -- wire
			Clock     : in  std_logic                    := 'X';             -- clk
			reset     : in  std_logic                    := 'X';             -- reset
			pixel_in  : in  std_logic_vector(7 downto 0) := (others => 'X'); -- wire
			eof_in    : in  std_logic                    := 'X';             -- wire
			sof_out   : out std_logic                                        -- wire
		);
	end component gaussian_ip_GN_gaussian_ip_Fusion_Decomposition_1;

	component gaussian_ip_GN_gaussian_ip_Fusion_Decomposition_2 is
		port (
			diff_in   : in  std_logic_vector(9 downto 0) := (others => 'X'); -- wire
			pixel_in  : in  std_logic_vector(7 downto 0) := (others => 'X'); -- wire
			eof_in    : in  std_logic                    := 'X';             -- wire
			sof_in    : in  std_logic                    := 'X';             -- wire
			diff_out  : out std_logic_vector(9 downto 0);                    -- wire
			valid_in  : in  std_logic                    := 'X';             -- wire
			valid_out : out std_logic;                                       -- wire
			sof_out   : out std_logic;                                       -- wire
			Clock     : in  std_logic                    := 'X';             -- clk
			reset     : in  std_logic                    := 'X';             -- reset
			eof_out   : out std_logic;                                       -- wire
			pixel_out : out std_logic_vector(7 downto 0)                     -- wire
		);
	end component gaussian_ip_GN_gaussian_ip_Fusion_Decomposition_2;

	component alt_dspbuilder_cast_GNBZR5PMEK is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(7 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(7 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNBZR5PMEK;

	component alt_dspbuilder_cast_GN46N4UJ5S is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic                    := 'X'; -- wire
			output : out std_logic_vector(0 downto 0)         -- wire
		);
	end component alt_dspbuilder_cast_GN46N4UJ5S;

	component alt_dspbuilder_cast_GN6DDKTPIR is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(7 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(9 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GN6DDKTPIR;

	signal multiplexeruser_aclrgnd_output_wire                 : std_logic;                    -- Multiplexeruser_aclrGND:output -> Multiplexer:user_aclr
	signal multiplexerenavcc_output_wire                       : std_logic;                    -- MultiplexerenaVCC:output -> Multiplexer:ena
	signal multiplexer1user_aclrgnd_output_wire                : std_logic;                    -- Multiplexer1user_aclrGND:output -> Multiplexer1:user_aclr
	signal multiplexer1enavcc_output_wire                      : std_logic;                    -- Multiplexer1enaVCC:output -> Multiplexer1:ena
	signal pipelined_adderuser_aclrgnd_output_wire             : std_logic;                    -- Pipelined_Adderuser_aclrGND:output -> Pipelined_Adder:user_aclr
	signal pipelined_adderenavcc_output_wire                   : std_logic;                    -- Pipelined_AdderenaVCC:output -> Pipelined_Adder:ena
	signal memory_delay3user_aclrgnd_output_wire               : std_logic;                    -- Memory_Delay3user_aclrGND:output -> Memory_Delay3:user_aclr
	signal memory_delay3enavcc_output_wire                     : std_logic;                    -- Memory_Delay3enaVCC:output -> Memory_Delay3:ena
	signal memory_delay1user_aclrgnd_output_wire               : std_logic;                    -- Memory_Delay1user_aclrGND:output -> Memory_Delay1:user_aclr
	signal memory_delay1enavcc_output_wire                     : std_logic;                    -- Memory_Delay1enaVCC:output -> Memory_Delay1:ena
	signal memory_delay2user_aclrgnd_output_wire               : std_logic;                    -- Memory_Delay2user_aclrGND:output -> Memory_Delay2:user_aclr
	signal memory_delay2enavcc_output_wire                     : std_logic;                    -- Memory_Delay2enaVCC:output -> Memory_Delay2:ena
	signal memory_delayuser_aclrgnd_output_wire                : std_logic;                    -- Memory_Delayuser_aclrGND:output -> Memory_Delay:user_aclr
	signal memory_delayenavcc_output_wire                      : std_logic;                    -- Memory_DelayenaVCC:output -> Memory_Delay:ena
	signal constant1_output_wire                               : std_logic_vector(9 downto 0); -- Constant1:output -> Comparator2:datab
	signal constant25_output_wire                              : std_logic_vector(1 downto 0); -- Constant25:output -> Bus_Concatenation1:a
	signal constant4_output_wire                               : std_logic_vector(9 downto 0); -- Constant4:output -> Comparator:datab
	signal gaussian_ip_fusion_decomposition_1_0_pixel_out_wire : std_logic_vector(7 downto 0); -- gaussian_ip_Fusion_Decomposition_1_0:pixel_out -> gaussian_ip_Fusion_Decomposition_2_0:pixel_in
	signal gaussian_ip_fusion_decomposition_1_0_diff_out_wire  : std_logic_vector(9 downto 0); -- gaussian_ip_Fusion_Decomposition_1_0:diff_out -> gaussian_ip_Fusion_Decomposition_2_0:diff_in
	signal gaussian_ip_fusion_decomposition_1_0_valid_out_wire : std_logic;                    -- gaussian_ip_Fusion_Decomposition_1_0:valid_out -> gaussian_ip_Fusion_Decomposition_2_0:valid_in
	signal gaussian_ip_fusion_decomposition_1_0_sof_out_wire   : std_logic;                    -- gaussian_ip_Fusion_Decomposition_1_0:sof_out -> gaussian_ip_Fusion_Decomposition_2_0:sof_in
	signal gaussian_ip_fusion_decomposition_1_0_eof_out_wire   : std_logic;                    -- gaussian_ip_Fusion_Decomposition_1_0:eof_out -> gaussian_ip_Fusion_Decomposition_2_0:eof_in
	signal gaussian_ip_fusion_decomposition_2_0_pixel_out_wire : std_logic_vector(7 downto 0); -- gaussian_ip_Fusion_Decomposition_2_0:pixel_out -> gaussian_ip_Fusion_Decomposition_3_0:pixel_in
	signal gaussian_ip_fusion_decomposition_2_0_diff_out_wire  : std_logic_vector(9 downto 0); -- gaussian_ip_Fusion_Decomposition_2_0:diff_out -> gaussian_ip_Fusion_Decomposition_3_0:diff_in
	signal gaussian_ip_fusion_decomposition_2_0_valid_out_wire : std_logic;                    -- gaussian_ip_Fusion_Decomposition_2_0:valid_out -> gaussian_ip_Fusion_Decomposition_3_0:valid_in
	signal gaussian_ip_fusion_decomposition_2_0_sof_out_wire   : std_logic;                    -- gaussian_ip_Fusion_Decomposition_2_0:sof_out -> gaussian_ip_Fusion_Decomposition_3_0:sof_in
	signal gaussian_ip_fusion_decomposition_2_0_eof_out_wire   : std_logic;                    -- gaussian_ip_Fusion_Decomposition_2_0:eof_out -> gaussian_ip_Fusion_Decomposition_3_0:eof_in
	signal pixel1_in_0_output_wire                             : std_logic_vector(7 downto 0); -- pixel1_in_0:output -> gaussian_ip_Fusion_Decomposition_1_0:pixel_in
	signal pipelined_adder_result_wire                         : std_logic_vector(9 downto 0); -- Pipelined_Adder:result -> [Comparator2:dataa, Comparator:dataa, Multiplexer1:in0]
	signal valid1_in_0_output_wire                             : std_logic;                    -- valid1_in_0:output -> gaussian_ip_Fusion_Decomposition_1_0:valid_in
	signal sof1_in_0_output_wire                               : std_logic;                    -- sof1_in_0:output -> gaussian_ip_Fusion_Decomposition_1_0:sof_in
	signal eof1_in_0_output_wire                               : std_logic;                    -- eof1_in_0:output -> gaussian_ip_Fusion_Decomposition_1_0:eof_in
	signal gaussian_ip_fusion_decomposition_3_0_diff_out_wire  : std_logic_vector(9 downto 0); -- gaussian_ip_Fusion_Decomposition_3_0:diff_out -> Memory_Delay:input
	signal multiplexer1_result_wire                            : std_logic_vector(9 downto 0); -- Multiplexer1:result -> Multiplexer:in0
	signal bus_concatenation1_output_wire                      : std_logic_vector(9 downto 0); -- Bus_Concatenation1:output -> Pipelined_Adder:dataa
	signal memory_delay_output_wire                            : std_logic_vector(9 downto 0); -- Memory_Delay:output -> Pipelined_Adder:datab
	signal multiplexer_result_wire                             : std_logic_vector(9 downto 0); -- Multiplexer:result -> pixel_out_0:input
	signal memory_delay1_output_wire                           : std_logic_vector(0 downto 0); -- Memory_Delay1:output -> valid_out_0:input
	signal memory_delay2_output_wire                           : std_logic_vector(0 downto 0); -- Memory_Delay2:output -> sof_out_0:input
	signal memory_delay3_output_wire                           : std_logic_vector(0 downto 0); -- Memory_Delay3:output -> eof_out_0:input
	signal gaussian_ip_fusion_decomposition_3_0_valid_out_wire : std_logic;                    -- gaussian_ip_Fusion_Decomposition_3_0:valid_out -> [cast200:input, ready2_in_0:input]
	signal pixel2_in_0_output_wire                             : std_logic_vector(7 downto 0); -- pixel2_in_0:output -> cast199:input
	signal cast199_output_wire                                 : std_logic_vector(7 downto 0); -- cast199:output -> Bus_Concatenation1:b
	signal cast200_output_wire                                 : std_logic_vector(0 downto 0); -- cast200:output -> Memory_Delay1:input
	signal gaussian_ip_fusion_decomposition_3_0_sof_out_wire   : std_logic;                    -- gaussian_ip_Fusion_Decomposition_3_0:sof_out -> cast201:input
	signal cast201_output_wire                                 : std_logic_vector(0 downto 0); -- cast201:output -> Memory_Delay2:input
	signal gaussian_ip_fusion_decomposition_3_0_eof_out_wire   : std_logic;                    -- gaussian_ip_Fusion_Decomposition_3_0:eof_out -> cast202:input
	signal cast202_output_wire                                 : std_logic_vector(0 downto 0); -- cast202:output -> Memory_Delay3:input
	signal comparator_result_wire                              : std_logic;                    -- Comparator:result -> cast203:input
	signal cast203_output_wire                                 : std_logic_vector(0 downto 0); -- cast203:output -> Multiplexer:sel
	signal constant3_output_wire                               : std_logic_vector(7 downto 0); -- Constant3:output -> cast204:input
	signal cast204_output_wire                                 : std_logic_vector(9 downto 0); -- cast204:output -> Multiplexer:in1
	signal comparator2_result_wire                             : std_logic;                    -- Comparator2:result -> cast205:input
	signal cast205_output_wire                                 : std_logic_vector(0 downto 0); -- cast205:output -> Multiplexer1:sel
	signal constant2_output_wire                               : std_logic_vector(7 downto 0); -- Constant2:output -> cast206:input
	signal cast206_output_wire                                 : std_logic_vector(9 downto 0); -- cast206:output -> Multiplexer1:in1
	signal clock_0_clock_output_clk                            : std_logic;                    -- Clock_0:clock_out -> [Bus_Concatenation1:clock, Comparator2:clock, Comparator:clock, Memory_Delay1:clock, Memory_Delay2:clock, Memory_Delay3:clock, Memory_Delay:clock, Multiplexer1:clock, Multiplexer:clock, Pipelined_Adder:clock, gaussian_ip_Fusion_Decomposition_1_0:Clock, gaussian_ip_Fusion_Decomposition_2_0:Clock, gaussian_ip_Fusion_Decomposition_3_0:Clock]
	signal clock_0_clock_output_reset                          : std_logic;                    -- Clock_0:aclr_out -> [Bus_Concatenation1:aclr, Comparator2:sclr, Comparator:sclr, Memory_Delay1:aclr, Memory_Delay2:aclr, Memory_Delay3:aclr, Memory_Delay:aclr, Multiplexer1:aclr, Multiplexer:aclr, Pipelined_Adder:aclr, gaussian_ip_Fusion_Decomposition_1_0:reset, gaussian_ip_Fusion_Decomposition_2_0:reset, gaussian_ip_Fusion_Decomposition_3_0:reset]

begin

	clock_0 : component alt_dspbuilder_clock_GNQFU4PUDH
		port map (
			clock_out => clock_0_clock_output_clk,   -- clock_output.clk
			aclr_out  => clock_0_clock_output_reset, --             .reset
			clock     => Clock,                      --        clock.clk
			aclr      => reset                       --             .reset
		);

	eof_out_0 : component alt_dspbuilder_port_GNXAOKDYKC
		port map (
			input  => memory_delay3_output_wire, --  input.wire
			output => eof_out                    -- output.wire
		);

	pixel2_in_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => pixel2_in,               --  input.wire
			output => pixel2_in_0_output_wire  -- output.wire
		);

	multiplexer : component alt_dspbuilder_multiplexer_GNWZZP2IFI
		generic map (
			number_inputs          => 2,
			pipeline               => 0,
			width                  => 10,
			HDLTYPE                => "STD_LOGIC_VECTOR",
			use_one_hot_select_bus => 0
		)
		port map (
			clock     => clock_0_clock_output_clk,            -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,          --           .reset
			sel       => cast203_output_wire,                 --        sel.wire
			result    => multiplexer_result_wire,             --     result.wire
			ena       => multiplexerenavcc_output_wire,       --        ena.wire
			user_aclr => multiplexeruser_aclrgnd_output_wire, --  user_aclr.wire
			in0       => multiplexer1_result_wire,            --        in0.wire
			in1       => cast204_output_wire                  --        in1.wire
		);

	multiplexeruser_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplexeruser_aclrgnd_output_wire  -- output.wire
		);

	multiplexerenavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => multiplexerenavcc_output_wire  -- output.wire
		);

	multiplexer1 : component alt_dspbuilder_multiplexer_GNWZZP2IFI
		generic map (
			number_inputs          => 2,
			pipeline               => 0,
			width                  => 10,
			HDLTYPE                => "STD_LOGIC_VECTOR",
			use_one_hot_select_bus => 0
		)
		port map (
			clock     => clock_0_clock_output_clk,             -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,           --           .reset
			sel       => cast205_output_wire,                  --        sel.wire
			result    => multiplexer1_result_wire,             --     result.wire
			ena       => multiplexer1enavcc_output_wire,       --        ena.wire
			user_aclr => multiplexer1user_aclrgnd_output_wire, --  user_aclr.wire
			in0       => pipelined_adder_result_wire,          --        in0.wire
			in1       => cast206_output_wire                   --        in1.wire
		);

	multiplexer1user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplexer1user_aclrgnd_output_wire  -- output.wire
		);

	multiplexer1enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => multiplexer1enavcc_output_wire  -- output.wire
		);

	ready2_in_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => gaussian_ip_fusion_decomposition_3_0_valid_out_wire, --  input.wire
			output => ready2_in                                            -- output.wire
		);

	constant25 : component alt_dspbuilder_constant_GN6SFEINY6
		generic map (
			BitPattern => "00",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 2
		)
		port map (
			output => constant25_output_wire  -- output.wire
		);

	pipelined_adder : component alt_dspbuilder_pipelined_adder_GN4HTUTWRG
		generic map (
			pipeline => 1,
			width    => 10
		)
		port map (
			clock     => clock_0_clock_output_clk,                -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,              --           .reset
			dataa     => bus_concatenation1_output_wire,          --      dataa.wire
			datab     => memory_delay_output_wire,                --      datab.wire
			result    => pipelined_adder_result_wire,             --     result.wire
			user_aclr => pipelined_adderuser_aclrgnd_output_wire, --  user_aclr.wire
			ena       => pipelined_adderenavcc_output_wire        --        ena.wire
		);

	pipelined_adderuser_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => pipelined_adderuser_aclrgnd_output_wire  -- output.wire
		);

	pipelined_adderenavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => pipelined_adderenavcc_output_wire  -- output.wire
		);

	comparator : component alt_dspbuilder_comparator_GN
		generic map (
			Operator  => "Altagb",
			lpm_width => 10
		)
		port map (
			clock  => clock_0_clock_output_clk,    -- clock_sclr.clk
			sclr   => clock_0_clock_output_reset,  --           .reset
			dataa  => pipelined_adder_result_wire, --      dataa.wire
			datab  => constant4_output_wire,       --      datab.wire
			result => comparator_result_wire       --     result.wire
		);

	valid_out_0 : component alt_dspbuilder_port_GNXAOKDYKC
		port map (
			input  => memory_delay1_output_wire, --  input.wire
			output => valid_out                  -- output.wire
		);

	memory_delay3 : component alt_dspbuilder_memdelay_GNR55NYJWV
		generic map (
			RAMTYPE => "AUTO",
			WIDTH   => 1,
			DELAY   => 2
		)
		port map (
			clock     => clock_0_clock_output_clk,              -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,            --           .reset
			input     => cast202_output_wire,                   --      input.wire
			output    => memory_delay3_output_wire,             --     output.wire
			user_aclr => memory_delay3user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => memory_delay3enavcc_output_wire        --        ena.wire
		);

	memory_delay3user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => memory_delay3user_aclrgnd_output_wire  -- output.wire
		);

	memory_delay3enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => memory_delay3enavcc_output_wire  -- output.wire
		);

	memory_delay1 : component alt_dspbuilder_memdelay_GNR55NYJWV
		generic map (
			RAMTYPE => "AUTO",
			WIDTH   => 1,
			DELAY   => 2
		)
		port map (
			clock     => clock_0_clock_output_clk,              -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,            --           .reset
			input     => cast200_output_wire,                   --      input.wire
			output    => memory_delay1_output_wire,             --     output.wire
			user_aclr => memory_delay1user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => memory_delay1enavcc_output_wire        --        ena.wire
		);

	memory_delay1user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => memory_delay1user_aclrgnd_output_wire  -- output.wire
		);

	memory_delay1enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => memory_delay1enavcc_output_wire  -- output.wire
		);

	comparator2 : component alt_dspbuilder_comparator_GN
		generic map (
			Operator  => "Altalb",
			lpm_width => 10
		)
		port map (
			clock  => clock_0_clock_output_clk,    -- clock_sclr.clk
			sclr   => clock_0_clock_output_reset,  --           .reset
			dataa  => pipelined_adder_result_wire, --      dataa.wire
			datab  => constant1_output_wire,       --      datab.wire
			result => comparator2_result_wire      --     result.wire
		);

	memory_delay2 : component alt_dspbuilder_memdelay_GNR55NYJWV
		generic map (
			RAMTYPE => "AUTO",
			WIDTH   => 1,
			DELAY   => 2
		)
		port map (
			clock     => clock_0_clock_output_clk,              -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,            --           .reset
			input     => cast201_output_wire,                   --      input.wire
			output    => memory_delay2_output_wire,             --     output.wire
			user_aclr => memory_delay2user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => memory_delay2enavcc_output_wire        --        ena.wire
		);

	memory_delay2user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => memory_delay2user_aclrgnd_output_wire  -- output.wire
		);

	memory_delay2enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => memory_delay2enavcc_output_wire  -- output.wire
		);

	eof1_in_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => eof1_in,               --  input.wire
			output => eof1_in_0_output_wire  -- output.wire
		);

	pixel1_in_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => pixel1_in,               --  input.wire
			output => pixel1_in_0_output_wire  -- output.wire
		);

	constant2 : component alt_dspbuilder_constant_GNC5NOVIJT
		generic map (
			BitPattern => "00000000",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 8
		)
		port map (
			output => constant2_output_wire  -- output.wire
		);

	constant3 : component alt_dspbuilder_constant_GNSVSRQZMI
		generic map (
			BitPattern => "11111111",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 8
		)
		port map (
			output => constant3_output_wire  -- output.wire
		);

	constant1 : component alt_dspbuilder_constant_GN5IRMZXKK
		generic map (
			BitPattern => "0000000000",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 10
		)
		port map (
			output => constant1_output_wire  -- output.wire
		);

	valid1_in_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => valid1_in,               --  input.wire
			output => valid1_in_0_output_wire  -- output.wire
		);

	bus_concatenation1 : component alt_dspbuilder_bus_concat_GNKLOJ6ING
		generic map (
			widthA => 2,
			widthB => 8
		)
		port map (
			clock  => clock_0_clock_output_clk,       -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,     --           .reset
			a      => constant25_output_wire,         --          a.wire
			b      => cast199_output_wire,            --          b.wire
			output => bus_concatenation1_output_wire  --     output.wire
		);

	sof1_in_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => sof1_in,               --  input.wire
			output => sof1_in_0_output_wire  -- output.wire
		);

	constant4 : component alt_dspbuilder_constant_GNK57PM5EK
		generic map (
			BitPattern => "0011111111",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 10
		)
		port map (
			output => constant4_output_wire  -- output.wire
		);

	memory_delay : component alt_dspbuilder_memdelay_GNT3M75IMA
		generic map (
			RAMTYPE => "AUTO",
			WIDTH   => 10,
			DELAY   => 1
		)
		port map (
			clock     => clock_0_clock_output_clk,                           -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,                         --           .reset
			input     => gaussian_ip_fusion_decomposition_3_0_diff_out_wire, --      input.wire
			output    => memory_delay_output_wire,                           --     output.wire
			user_aclr => memory_delayuser_aclrgnd_output_wire,               --  user_aclr.wire
			ena       => memory_delayenavcc_output_wire                      --        ena.wire
		);

	memory_delayuser_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => memory_delayuser_aclrgnd_output_wire  -- output.wire
		);

	memory_delayenavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => memory_delayenavcc_output_wire  -- output.wire
		);

	sof_out_0 : component alt_dspbuilder_port_GNXAOKDYKC
		port map (
			input  => memory_delay2_output_wire, --  input.wire
			output => sof_out                    -- output.wire
		);

	pixel_out_0 : component alt_dspbuilder_port_GNSSYS4J5R
		port map (
			input  => multiplexer_result_wire, --  input.wire
			output => pixel_out                -- output.wire
		);

	gaussian_ip_fusion_decomposition_3_0 : component gaussian_ip_GN_gaussian_ip_Fusion_Decomposition_3
		port map (
			sof_in    => gaussian_ip_fusion_decomposition_2_0_sof_out_wire,   --    sof_in.wire
			sof_out   => gaussian_ip_fusion_decomposition_3_0_sof_out_wire,   --   sof_out.wire
			Clock     => clock_0_clock_output_clk,                            --     Clock.clk
			reset     => clock_0_clock_output_reset,                          --          .reset
			eof_in    => gaussian_ip_fusion_decomposition_2_0_eof_out_wire,   --    eof_in.wire
			eof_out   => gaussian_ip_fusion_decomposition_3_0_eof_out_wire,   --   eof_out.wire
			valid_in  => gaussian_ip_fusion_decomposition_2_0_valid_out_wire, --  valid_in.wire
			diff_out  => gaussian_ip_fusion_decomposition_3_0_diff_out_wire,  --  diff_out.wire
			valid_out => gaussian_ip_fusion_decomposition_3_0_valid_out_wire, -- valid_out.wire
			diff_in   => gaussian_ip_fusion_decomposition_2_0_diff_out_wire,  --   diff_in.wire
			pixel_out => open,                                                -- pixel_out.wire
			pixel_in  => gaussian_ip_fusion_decomposition_2_0_pixel_out_wire  --  pixel_in.wire
		);

	gaussian_ip_fusion_decomposition_1_0 : component gaussian_ip_GN_gaussian_ip_Fusion_Decomposition_1
		port map (
			valid_in  => valid1_in_0_output_wire,                             --  valid_in.wire
			valid_out => gaussian_ip_fusion_decomposition_1_0_valid_out_wire, -- valid_out.wire
			pixel_out => gaussian_ip_fusion_decomposition_1_0_pixel_out_wire, -- pixel_out.wire
			diff_out  => gaussian_ip_fusion_decomposition_1_0_diff_out_wire,  --  diff_out.wire
			eof_out   => gaussian_ip_fusion_decomposition_1_0_eof_out_wire,   --   eof_out.wire
			sof_in    => sof1_in_0_output_wire,                               --    sof_in.wire
			Clock     => clock_0_clock_output_clk,                            --     Clock.clk
			reset     => clock_0_clock_output_reset,                          --          .reset
			pixel_in  => pixel1_in_0_output_wire,                             --  pixel_in.wire
			eof_in    => eof1_in_0_output_wire,                               --    eof_in.wire
			sof_out   => gaussian_ip_fusion_decomposition_1_0_sof_out_wire    --   sof_out.wire
		);

	gaussian_ip_fusion_decomposition_2_0 : component gaussian_ip_GN_gaussian_ip_Fusion_Decomposition_2
		port map (
			diff_in   => gaussian_ip_fusion_decomposition_1_0_diff_out_wire,  --   diff_in.wire
			pixel_in  => gaussian_ip_fusion_decomposition_1_0_pixel_out_wire, --  pixel_in.wire
			eof_in    => gaussian_ip_fusion_decomposition_1_0_eof_out_wire,   --    eof_in.wire
			sof_in    => gaussian_ip_fusion_decomposition_1_0_sof_out_wire,   --    sof_in.wire
			diff_out  => gaussian_ip_fusion_decomposition_2_0_diff_out_wire,  --  diff_out.wire
			valid_in  => gaussian_ip_fusion_decomposition_1_0_valid_out_wire, --  valid_in.wire
			valid_out => gaussian_ip_fusion_decomposition_2_0_valid_out_wire, -- valid_out.wire
			sof_out   => gaussian_ip_fusion_decomposition_2_0_sof_out_wire,   --   sof_out.wire
			Clock     => clock_0_clock_output_clk,                            --     Clock.clk
			reset     => clock_0_clock_output_reset,                          --          .reset
			eof_out   => gaussian_ip_fusion_decomposition_2_0_eof_out_wire,   --   eof_out.wire
			pixel_out => gaussian_ip_fusion_decomposition_2_0_pixel_out_wire  -- pixel_out.wire
		);

	cast199 : component alt_dspbuilder_cast_GNBZR5PMEK
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => pixel2_in_0_output_wire, --  input.wire
			output => cast199_output_wire      -- output.wire
		);

	cast200 : component alt_dspbuilder_cast_GN46N4UJ5S
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => gaussian_ip_fusion_decomposition_3_0_valid_out_wire, --  input.wire
			output => cast200_output_wire                                  -- output.wire
		);

	cast201 : component alt_dspbuilder_cast_GN46N4UJ5S
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => gaussian_ip_fusion_decomposition_3_0_sof_out_wire, --  input.wire
			output => cast201_output_wire                                -- output.wire
		);

	cast202 : component alt_dspbuilder_cast_GN46N4UJ5S
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => gaussian_ip_fusion_decomposition_3_0_eof_out_wire, --  input.wire
			output => cast202_output_wire                                -- output.wire
		);

	cast203 : component alt_dspbuilder_cast_GN46N4UJ5S
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => comparator_result_wire, --  input.wire
			output => cast203_output_wire     -- output.wire
		);

	cast204 : component alt_dspbuilder_cast_GN6DDKTPIR
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => constant3_output_wire, --  input.wire
			output => cast204_output_wire    -- output.wire
		);

	cast205 : component alt_dspbuilder_cast_GN46N4UJ5S
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => comparator2_result_wire, --  input.wire
			output => cast205_output_wire      -- output.wire
		);

	cast206 : component alt_dspbuilder_cast_GN6DDKTPIR
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => constant2_output_wire, --  input.wire
			output => cast206_output_wire    -- output.wire
		);

end architecture rtl; -- of gaussian_ip_GN_gaussian_ip_Fusion
