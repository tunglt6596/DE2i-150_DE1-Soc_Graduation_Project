-- localedgepreserve_GN_localedgepreserve_Fusion_Cal_A_B_2.vhd

-- Generated using ACDS version 17.1 590

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity localedgepreserve_GN_localedgepreserve_Fusion_Cal_A_B_2 is
	port (
		eof_in    : in  std_logic                     := '0';             --    eof_in.wire
		a_out     : out std_logic_vector(15 downto 0);                    --     a_out.wire
		pixel_in  : in  std_logic_vector(7 downto 0)  := (others => '0'); --  pixel_in.wire
		b_out     : out std_logic_vector(15 downto 0);                    --     b_out.wire
		pixel_out : out std_logic_vector(7 downto 0);                     -- pixel_out.wire
		Clock     : in  std_logic                     := '0';             --     Clock.clk
		reset     : in  std_logic                     := '0';             --          .reset
		grad_in   : in  std_logic_vector(10 downto 0) := (others => '0'); --   grad_in.wire
		eof_out   : out std_logic;                                        --   eof_out.wire
		valid_in  : in  std_logic                     := '0';             --  valid_in.wire
		valid_out : out std_logic                                         -- valid_out.wire
	);
end entity localedgepreserve_GN_localedgepreserve_Fusion_Cal_A_B_2;

architecture rtl of localedgepreserve_GN_localedgepreserve_Fusion_Cal_A_B_2 is
	component alt_dspbuilder_clock_GNQFU4PUDH is
		port (
			aclr      : in  std_logic := 'X'; -- reset
			aclr_n    : in  std_logic := 'X'; -- reset_n
			aclr_out  : out std_logic;        -- reset
			clock     : in  std_logic := 'X'; -- clk
			clock_out : out std_logic         -- clk
		);
	end component alt_dspbuilder_clock_GNQFU4PUDH;

	component alt_dspbuilder_port_GN37ALZBS4 is
		port (
			input  : in  std_logic := 'X'; -- wire
			output : out std_logic         -- wire
		);
	end component alt_dspbuilder_port_GN37ALZBS4;

	component alt_dspbuilder_multiplier_GN2GJCFTFE is
		generic (
			aWidth                         : natural := 8;
			Signed                         : natural := 0;
			bWidth                         : natural := 8;
			DEDICATED_MULTIPLIER_CIRCUITRY : string  := "AUTO";
			pipeline                       : integer := 0;
			OutputLsb                      : integer := 0;
			OutputMsb                      : integer := 8
		);
		port (
			aclr      : in  std_logic                                          := 'X';             -- clk
			clock     : in  std_logic                                          := 'X';             -- clk
			dataa     : in  std_logic_vector(aWidth-1 downto 0)                := (others => 'X'); -- wire
			datab     : in  std_logic_vector(bWidth-1 downto 0)                := (others => 'X'); -- wire
			ena       : in  std_logic                                          := 'X';             -- wire
			result    : out std_logic_vector(OutputMsb-OutputLsb+1-1 downto 0);                    -- wire
			user_aclr : in  std_logic                                          := 'X'              -- wire
		);
	end component alt_dspbuilder_multiplier_GN2GJCFTFE;

	component alt_dspbuilder_gnd_GN is
		port (
			output : out std_logic   -- wire
		);
	end component alt_dspbuilder_gnd_GN;

	component alt_dspbuilder_cast_GNUYRTQ4QH is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(23 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNUYRTQ4QH;

	component alt_dspbuilder_multiplexer_GN7X7SG76C is
		generic (
			number_inputs          : natural  := 4;
			pipeline               : natural  := 0;
			width                  : positive := 8;
			HDLTYPE                : string   := "STD_LOGIC_VECTOR";
			use_one_hot_select_bus : natural  := 0
		);
		port (
			clock     : in  std_logic                     := 'X';             -- clk
			aclr      : in  std_logic                     := 'X';             -- reset
			sel       : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- wire
			result    : out std_logic_vector(15 downto 0);                    -- wire
			ena       : in  std_logic                     := 'X';             -- wire
			user_aclr : in  std_logic                     := 'X';             -- wire
			in0       : in  std_logic_vector(15 downto 0) := (others => 'X'); -- wire
			in1       : in  std_logic_vector(15 downto 0) := (others => 'X')  -- wire
		);
	end component alt_dspbuilder_multiplexer_GN7X7SG76C;

	component alt_dspbuilder_vcc_GN is
		port (
			output : out std_logic   -- wire
		);
	end component alt_dspbuilder_vcc_GN;

	component alt_dspbuilder_port_GNLA26EJAH is
		port (
			input  : in  std_logic_vector(10 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(10 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNLA26EJAH;

	component alt_dspbuilder_port_GNA5S4SQDN is
		port (
			input  : in  std_logic_vector(7 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(7 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNA5S4SQDN;

	component alt_dspbuilder_memdelay_GNDI52L3LZ is
		generic (
			RAMTYPE : string   := "AUTO";
			WIDTH   : positive := 8;
			DELAY   : positive := 1
		);
		port (
			aclr      : in  std_logic                          := 'X';             -- clk
			clock     : in  std_logic                          := 'X';             -- clk
			ena       : in  std_logic                          := 'X';             -- wire
			input     : in  std_logic_vector(WIDTH-1 downto 0) := (others => 'X'); -- wire
			output    : out std_logic_vector(WIDTH-1 downto 0);                    -- wire
			user_aclr : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_memdelay_GNDI52L3LZ;

	component alt_dspbuilder_pipelined_adder_GNTWZRTG4I is
		generic (
			pipeline : integer := 0;
			width    : natural := 0
		);
		port (
			aclr      : in  std_logic                          := 'X';             -- clk
			add_sub   : in  std_logic                          := 'X';             -- wire
			cin       : in  std_logic                          := 'X';             -- wire
			clock     : in  std_logic                          := 'X';             -- clk
			cout      : out std_logic;                                             -- wire
			dataa     : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			datab     : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			ena       : in  std_logic                          := 'X';             -- wire
			result    : out std_logic_vector(width-1 downto 0);                    -- wire
			user_aclr : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_pipelined_adder_GNTWZRTG4I;

	component alt_dspbuilder_memdelay_GNMIZKWFE6 is
		generic (
			RAMTYPE : string   := "AUTO";
			WIDTH   : positive := 8;
			DELAY   : positive := 1
		);
		port (
			aclr      : in  std_logic                          := 'X';             -- clk
			clock     : in  std_logic                          := 'X';             -- clk
			ena       : in  std_logic                          := 'X';             -- wire
			input     : in  std_logic_vector(WIDTH-1 downto 0) := (others => 'X'); -- wire
			output    : out std_logic_vector(WIDTH-1 downto 0);                    -- wire
			user_aclr : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_memdelay_GNMIZKWFE6;

	component alt_dspbuilder_memdelay_GNI6WYI4F7 is
		generic (
			RAMTYPE : string   := "AUTO";
			WIDTH   : positive := 8;
			DELAY   : positive := 1
		);
		port (
			aclr      : in  std_logic                          := 'X';             -- clk
			clock     : in  std_logic                          := 'X';             -- clk
			ena       : in  std_logic                          := 'X';             -- wire
			input     : in  std_logic_vector(WIDTH-1 downto 0) := (others => 'X'); -- wire
			output    : out std_logic_vector(WIDTH-1 downto 0);                    -- wire
			user_aclr : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_memdelay_GNI6WYI4F7;

	component localedgepreserve_GN_localedgepreserve_Fusion_Cal_A_B_2_Cal_MeanI_VarI is
		port (
			valid_in  : in  std_logic                     := 'X';             -- wire
			Clock     : in  std_logic                     := 'X';             -- clk
			reset     : in  std_logic                     := 'X';             -- reset
			pixel_out : out std_logic_vector(7 downto 0);                     -- wire
			pixel_in  : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- wire
			varI      : out std_logic_vector(39 downto 0);                    -- wire
			meanI     : out std_logic_vector(31 downto 0)                     -- wire
		);
	end component localedgepreserve_GN_localedgepreserve_Fusion_Cal_A_B_2_Cal_MeanI_VarI;

	component alt_dspbuilder_memdelay_GNF7HJJOOI is
		generic (
			RAMTYPE : string   := "AUTO";
			WIDTH   : positive := 8;
			DELAY   : positive := 1
		);
		port (
			aclr      : in  std_logic                          := 'X';             -- clk
			clock     : in  std_logic                          := 'X';             -- clk
			ena       : in  std_logic                          := 'X';             -- wire
			input     : in  std_logic_vector(WIDTH-1 downto 0) := (others => 'X'); -- wire
			output    : out std_logic_vector(WIDTH-1 downto 0);                    -- wire
			user_aclr : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_memdelay_GNF7HJJOOI;

	component alt_dspbuilder_comparator_GN is
		generic (
			Operator  : string  := "Altaeb";
			lpm_width : natural := 8
		);
		port (
			clock  : in  std_logic                              := 'X';             -- clk
			dataa  : in  std_logic_vector(lpm_width-1 downto 0) := (others => 'X'); -- wire
			datab  : in  std_logic_vector(lpm_width-1 downto 0) := (others => 'X'); -- wire
			result : out std_logic;                                                 -- wire
			sclr   : in  std_logic                              := 'X'              -- clk
		);
	end component alt_dspbuilder_comparator_GN;

	component alt_dspbuilder_memdelay_GN4TPDAUQN is
		generic (
			RAMTYPE : string   := "AUTO";
			WIDTH   : positive := 8;
			DELAY   : positive := 1
		);
		port (
			aclr      : in  std_logic                          := 'X';             -- clk
			clock     : in  std_logic                          := 'X';             -- clk
			ena       : in  std_logic                          := 'X';             -- wire
			input     : in  std_logic_vector(WIDTH-1 downto 0) := (others => 'X'); -- wire
			output    : out std_logic_vector(WIDTH-1 downto 0);                    -- wire
			user_aclr : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_memdelay_GN4TPDAUQN;

	component alt_dspbuilder_memdelay_GNMYXI7BAD is
		generic (
			RAMTYPE : string   := "AUTO";
			WIDTH   : positive := 8;
			DELAY   : positive := 1
		);
		port (
			aclr      : in  std_logic                          := 'X';             -- clk
			clock     : in  std_logic                          := 'X';             -- clk
			ena       : in  std_logic                          := 'X';             -- wire
			input     : in  std_logic_vector(WIDTH-1 downto 0) := (others => 'X'); -- wire
			output    : out std_logic_vector(WIDTH-1 downto 0);                    -- wire
			user_aclr : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_memdelay_GNMYXI7BAD;

	component alt_dspbuilder_memdelay_GNNY7HWC5A is
		generic (
			RAMTYPE : string   := "AUTO";
			WIDTH   : positive := 8;
			DELAY   : positive := 1
		);
		port (
			aclr      : in  std_logic                          := 'X';             -- clk
			clock     : in  std_logic                          := 'X';             -- clk
			ena       : in  std_logic                          := 'X';             -- wire
			input     : in  std_logic_vector(WIDTH-1 downto 0) := (others => 'X'); -- wire
			output    : out std_logic_vector(WIDTH-1 downto 0);                    -- wire
			user_aclr : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_memdelay_GNNY7HWC5A;

	component alt_dspbuilder_memdelay_GNZWVQQT43 is
		generic (
			RAMTYPE : string   := "AUTO";
			WIDTH   : positive := 8;
			DELAY   : positive := 1
		);
		port (
			aclr      : in  std_logic                          := 'X';             -- clk
			clock     : in  std_logic                          := 'X';             -- clk
			ena       : in  std_logic                          := 'X';             -- wire
			input     : in  std_logic_vector(WIDTH-1 downto 0) := (others => 'X'); -- wire
			output    : out std_logic_vector(WIDTH-1 downto 0);                    -- wire
			user_aclr : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_memdelay_GNZWVQQT43;

	component alt_dspbuilder_multiplier_GNKTEWW72G is
		generic (
			aWidth                         : natural := 8;
			Signed                         : natural := 0;
			bWidth                         : natural := 8;
			DEDICATED_MULTIPLIER_CIRCUITRY : string  := "AUTO";
			pipeline                       : integer := 0;
			OutputLsb                      : integer := 0;
			OutputMsb                      : integer := 8
		);
		port (
			aclr      : in  std_logic                                          := 'X';             -- clk
			clock     : in  std_logic                                          := 'X';             -- clk
			dataa     : in  std_logic_vector(aWidth-1 downto 0)                := (others => 'X'); -- wire
			datab     : in  std_logic_vector(bWidth-1 downto 0)                := (others => 'X'); -- wire
			ena       : in  std_logic                                          := 'X';             -- wire
			result    : out std_logic_vector(OutputMsb-OutputLsb+1-1 downto 0);                    -- wire
			user_aclr : in  std_logic                                          := 'X'              -- wire
		);
	end component alt_dspbuilder_multiplier_GNKTEWW72G;

	component alt_dspbuilder_pipelined_adder_GNWEIMU3MK is
		generic (
			pipeline : integer := 0;
			width    : natural := 0
		);
		port (
			aclr      : in  std_logic                          := 'X';             -- clk
			add_sub   : in  std_logic                          := 'X';             -- wire
			cin       : in  std_logic                          := 'X';             -- wire
			clock     : in  std_logic                          := 'X';             -- clk
			cout      : out std_logic;                                             -- wire
			dataa     : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			datab     : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			ena       : in  std_logic                          := 'X';             -- wire
			result    : out std_logic_vector(width-1 downto 0);                    -- wire
			user_aclr : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_pipelined_adder_GNWEIMU3MK;

	component alt_dspbuilder_cast_GNPPZDVXTY is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(15 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNPPZDVXTY;

	component alt_dspbuilder_cast_GNW6I55EUT is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(7 downto 0)                      -- wire
		);
	end component alt_dspbuilder_cast_GNW6I55EUT;

	component alt_dspbuilder_port_GNBO6OMO5Y is
		port (
			input  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(15 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNBO6OMO5Y;

	component alt_dspbuilder_cast_GNZYD62DLY is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(39 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(23 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNZYD62DLY;

	component localedgepreserve_GN_localedgepreserve_Fusion_Cal_A_B_2_Cal_MeanG is
		port (
			meanG    : out std_logic_vector(34 downto 0);                    -- wire
			Clock    : in  std_logic                     := 'X';             -- clk
			reset    : in  std_logic                     := 'X';             -- reset
			valid_in : in  std_logic                     := 'X';             -- wire
			pixel_in : in  std_logic_vector(10 downto 0) := (others => 'X')  -- wire
		);
	end component localedgepreserve_GN_localedgepreserve_Fusion_Cal_A_B_2_Cal_MeanG;

	component alt_dspbuilder_constant_GNRSDUIWRP is
		generic (
			BitPattern : string  := "0000";
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(31 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GNRSDUIWRP;

	component localedgepreserve_GN_localedgepreserve_Fusion_Cal_A_B_2_generate_signals is
		port (
			Clock     : in  std_logic := 'X'; -- clk
			reset     : in  std_logic := 'X'; -- reset
			valid_in  : in  std_logic := 'X'; -- wire
			eof_out   : out std_logic;        -- wire
			valid_out : out std_logic;        -- wire
			eof_in    : in  std_logic := 'X'  -- wire
		);
	end component localedgepreserve_GN_localedgepreserve_Fusion_Cal_A_B_2_generate_signals;

	component alt_dspbuilder_bus_concat_GNOQTN4QAD is
		generic (
			widthA : natural := 8;
			widthB : natural := 8
		);
		port (
			a      : in  std_logic_vector(widthA-1 downto 0)        := (others => 'X'); -- wire
			aclr   : in  std_logic                                  := 'X';             -- clk
			b      : in  std_logic_vector(widthB-1 downto 0)        := (others => 'X'); -- wire
			clock  : in  std_logic                                  := 'X';             -- clk
			output : out std_logic_vector(widthA+widthB-1 downto 0)                     -- wire
		);
	end component alt_dspbuilder_bus_concat_GNOQTN4QAD;

	component alt_dspbuilder_bus_concat_GNDDREGCTK is
		generic (
			widthA : natural := 8;
			widthB : natural := 8
		);
		port (
			a      : in  std_logic_vector(widthA-1 downto 0)        := (others => 'X'); -- wire
			aclr   : in  std_logic                                  := 'X';             -- clk
			b      : in  std_logic_vector(widthB-1 downto 0)        := (others => 'X'); -- wire
			clock  : in  std_logic                                  := 'X';             -- clk
			output : out std_logic_vector(widthA+widthB-1 downto 0)                     -- wire
		);
	end component alt_dspbuilder_bus_concat_GNDDREGCTK;

	component alt_dspbuilder_constant_GNC5NOVIJT is
		generic (
			BitPattern : string  := "0000";
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(7 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GNC5NOVIJT;

	component alt_dspbuilder_constant_GNCWI5QDAD is
		generic (
			BitPattern : string  := "0000";
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(15 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GNCWI5QDAD;

	component alt_dspbuilder_constant_GN5FET4EJH is
		generic (
			BitPattern : string  := "0000";
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(23 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GN5FET4EJH;

	component div is
		port (
			clk : in  std_logic                     := 'X';             -- clk
			d   : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			ena : in  std_logic                     := 'X';             -- wire
			q   : out std_logic_vector(23 downto 0);                    -- wire
			z   : in  std_logic_vector(47 downto 0) := (others => 'X')  -- wire
		);
	end component div;

	component alt_dspbuilder_cast_GN3FODBL3U is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(40 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GN3FODBL3U;

	component alt_dspbuilder_cast_GNKD3JEUSD is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(47 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(47 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNKD3JEUSD;

	component alt_dspbuilder_cast_GN5P6ORZXA is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(23 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GN5P6ORZXA;

	component alt_dspbuilder_cast_GNEIIG67TZ is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(23 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNEIIG67TZ;

	component alt_dspbuilder_cast_GNOEMJJSIT is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(39 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(39 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNOEMJJSIT;

	component alt_dspbuilder_cast_GNA5TAMWCZ is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(23 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNA5TAMWCZ;

	component alt_dspbuilder_cast_GNP5J2CFQQ is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(40 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNP5J2CFQQ;

	component alt_dspbuilder_cast_GN46N4UJ5S is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic                    := 'X'; -- wire
			output : out std_logic_vector(0 downto 0)         -- wire
		);
	end component alt_dspbuilder_cast_GN46N4UJ5S;

	component alt_dspbuilder_cast_GNDHESB5KA is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- wire
			output : out std_logic_vector(15 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNDHESB5KA;

	component alt_dspbuilder_cast_GNT7Y2ULVV is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(7 downto 0)                      -- wire
		);
	end component alt_dspbuilder_cast_GNT7Y2ULVV;

	component alt_dspbuilder_cast_GNXSA7APAK is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(34 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(39 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNXSA7APAK;

	signal multiplier1user_aclrgnd_output_wire                                  : std_logic;                     -- Multiplier1user_aclrGND:output -> Multiplier1:user_aclr
	signal multiplexeruser_aclrgnd_output_wire                                  : std_logic;                     -- Multiplexeruser_aclrGND:output -> Multiplexer:user_aclr
	signal multiplexerenavcc_output_wire                                        : std_logic;                     -- MultiplexerenaVCC:output -> Multiplexer:ena
	signal memory_delay7user_aclrgnd_output_wire                                : std_logic;                     -- Memory_Delay7user_aclrGND:output -> Memory_Delay7:user_aclr
	signal pipelined_adderuser_aclrgnd_output_wire                              : std_logic;                     -- Pipelined_Adderuser_aclrGND:output -> Pipelined_Adder:user_aclr
	signal memory_delay5user_aclrgnd_output_wire                                : std_logic;                     -- Memory_Delay5user_aclrGND:output -> Memory_Delay5:user_aclr
	signal memory_delay6user_aclrgnd_output_wire                                : std_logic;                     -- Memory_Delay6user_aclrGND:output -> Memory_Delay6:user_aclr
	signal memory_delay9user_aclrgnd_output_wire                                : std_logic;                     -- Memory_Delay9user_aclrGND:output -> Memory_Delay9:user_aclr
	signal memory_delay3user_aclrgnd_output_wire                                : std_logic;                     -- Memory_Delay3user_aclrGND:output -> Memory_Delay3:user_aclr
	signal memory_delay4user_aclrgnd_output_wire                                : std_logic;                     -- Memory_Delay4user_aclrGND:output -> Memory_Delay4:user_aclr
	signal memory_delay1user_aclrgnd_output_wire                                : std_logic;                     -- Memory_Delay1user_aclrGND:output -> Memory_Delay1:user_aclr
	signal memory_delay2user_aclrgnd_output_wire                                : std_logic;                     -- Memory_Delay2user_aclrGND:output -> Memory_Delay2:user_aclr
	signal multiplieruser_aclrgnd_output_wire                                   : std_logic;                     -- Multiplieruser_aclrGND:output -> Multiplier:user_aclr
	signal pipelined_adder1user_aclrgnd_output_wire                             : std_logic;                     -- Pipelined_Adder1user_aclrGND:output -> Pipelined_Adder1:user_aclr
	signal bus_concatenation2_output_wire                                       : std_logic_vector(31 downto 0); -- Bus_Concatenation2:output -> Bus_Concatenation3:b
	signal bus_conversion2_output_wire                                          : std_logic_vector(23 downto 0); -- Bus_Conversion2:output -> Binary_Point_Casting3:input
	signal bus_conversion3_output_wire                                          : std_logic_vector(23 downto 0); -- Bus_Conversion3:output -> Binary_Point_Casting2:input
	signal binary_point_casting1_output_wire                                    : std_logic_vector(23 downto 0); -- Binary_Point_Casting1:output -> Bus_Conversion4:input
	signal constant6_output_wire                                                : std_logic_vector(7 downto 0);  -- Constant6:output -> Bus_Concatenation2:b
	signal constant7_output_wire                                                : std_logic_vector(15 downto 0); -- Constant7:output -> Bus_Concatenation3:a
	signal grad_in_0_output_wire                                                : std_logic_vector(10 downto 0); -- grad_in_0:output -> localedgepreserve_Fusion_Cal_A_B_2_Cal_MeanG_0:pixel_in
	signal localedgepreserve_fusion_cal_a_b_2_cal_meani_vari_0_meani_wire       : std_logic_vector(31 downto 0); -- localedgepreserve_Fusion_Cal_A_B_2_Cal_MeanI_VarI_0:meanI -> Bus_Conversion5:input
	signal valid_in_0_output_wire                                               : std_logic;                     -- valid_in_0:output -> [Divider:ena, Memory_Delay1:ena, Memory_Delay2:ena, Memory_Delay3:ena, Memory_Delay4:ena, Memory_Delay5:ena, Memory_Delay6:ena, Memory_Delay7:ena, Memory_Delay9:ena, Multiplier1:ena, Multiplier:ena, Pipelined_Adder1:ena, Pipelined_Adder:ena, localedgepreserve_Fusion_Cal_A_B_2_Cal_MeanG_0:valid_in, localedgepreserve_Fusion_Cal_A_B_2_Cal_MeanI_VarI_0:valid_in, localedgepreserve_Fusion_Cal_A_B_2_generate_signals_0:valid_in]
	signal pixel_in_0_output_wire                                               : std_logic_vector(7 downto 0);  -- pixel_in_0:output -> localedgepreserve_Fusion_Cal_A_B_2_Cal_MeanI_VarI_0:pixel_in
	signal localedgepreserve_fusion_cal_a_b_2_cal_meani_vari_0_vari_wire        : std_logic_vector(39 downto 0); -- localedgepreserve_Fusion_Cal_A_B_2_Cal_MeanI_VarI_0:varI -> Memory_Delay1:input
	signal binary_point_casting3_output_wire                                    : std_logic_vector(23 downto 0); -- Binary_Point_Casting3:output -> Memory_Delay2:input
	signal bus_conversion5_output_wire                                          : std_logic_vector(15 downto 0); -- Bus_Conversion5:output -> Memory_Delay3:input
	signal multiplexer_result_wire                                              : std_logic_vector(15 downto 0); -- Multiplexer:result -> [Memory_Delay4:input, cast115:input]
	signal memory_delay3_output_wire                                            : std_logic_vector(15 downto 0); -- Memory_Delay3:output -> [Memory_Delay5:input, Multiplier:dataa]
	signal localedgepreserve_fusion_cal_a_b_2_cal_meani_vari_0_pixel_out_wire   : std_logic_vector(7 downto 0);  -- localedgepreserve_Fusion_Cal_A_B_2_Cal_MeanI_VarI_0:pixel_out -> Memory_Delay6:input
	signal memory_delay2_output_wire                                            : std_logic_vector(23 downto 0); -- Memory_Delay2:output -> [Memory_Delay7:input, cast111:input]
	signal localedgepreserve_fusion_cal_a_b_2_cal_meang_0_meang_wire            : std_logic_vector(34 downto 0); -- localedgepreserve_Fusion_Cal_A_B_2_Cal_MeanG_0:meanG -> Memory_Delay9:input
	signal constant4_output_wire                                                : std_logic_vector(15 downto 0); -- Constant4:output -> Multiplexer:in1
	signal memory_delay9_output_wire                                            : std_logic_vector(34 downto 0); -- Memory_Delay9:output -> Multiplier1:dataa
	signal constant_1_output_wire                                               : std_logic_vector(23 downto 0); -- Constant_1:output -> Multiplier1:datab
	signal pipelined_adder_result_wire                                          : std_logic_vector(39 downto 0); -- Pipelined_Adder:result -> Bus_Conversion3:input
	signal memory_delay5_output_wire                                            : std_logic_vector(15 downto 0); -- Memory_Delay5:output -> Pipelined_Adder1:dataa
	signal multiplier_result_wire                                               : std_logic_vector(15 downto 0); -- Multiplier:result -> Pipelined_Adder1:datab
	signal eof_in_0_output_wire                                                 : std_logic;                     -- eof_in_0:output -> localedgepreserve_Fusion_Cal_A_B_2_generate_signals_0:eof_in
	signal memory_delay6_output_wire                                            : std_logic_vector(7 downto 0);  -- Memory_Delay6:output -> pixel_out_0:input
	signal memory_delay4_output_wire                                            : std_logic_vector(15 downto 0); -- Memory_Delay4:output -> a_out_0:input
	signal pipelined_adder1_result_wire                                         : std_logic_vector(15 downto 0); -- Pipelined_Adder1:result -> b_out_0:input
	signal localedgepreserve_fusion_cal_a_b_2_generate_signals_0_valid_out_wire : std_logic;                     -- localedgepreserve_Fusion_Cal_A_B_2_generate_signals_0:valid_out -> valid_out_0:input
	signal localedgepreserve_fusion_cal_a_b_2_generate_signals_0_eof_out_wire   : std_logic;                     -- localedgepreserve_Fusion_Cal_A_B_2_generate_signals_0:eof_out -> eof_out_0:input
	signal constant1_output_wire                                                : std_logic_vector(31 downto 0); -- Constant1:output -> cast106:input
	signal cast106_output_wire                                                  : std_logic_vector(40 downto 0); -- cast106:output -> Comparator:datab
	signal bus_concatenation3_output_wire                                       : std_logic_vector(47 downto 0); -- Bus_Concatenation3:output -> cast107:input
	signal cast107_output_wire                                                  : std_logic_vector(47 downto 0); -- cast107:output -> Divider:z
	signal binary_point_casting2_output_wire                                    : std_logic_vector(23 downto 0); -- Binary_Point_Casting2:output -> cast108:input
	signal cast108_output_wire                                                  : std_logic_vector(23 downto 0); -- cast108:output -> Divider:d
	signal divider_q_wire                                                       : std_logic_vector(23 downto 0); -- Divider:q -> cast109:input
	signal cast109_output_wire                                                  : std_logic_vector(23 downto 0); -- cast109:output -> Binary_Point_Casting1:input
	signal memory_delay1_output_wire                                            : std_logic_vector(39 downto 0); -- Memory_Delay1:output -> [cast110:input, cast116:input]
	signal cast110_output_wire                                                  : std_logic_vector(39 downto 0); -- cast110:output -> Bus_Conversion2:input
	signal cast111_output_wire                                                  : std_logic_vector(23 downto 0); -- cast111:output -> Bus_Concatenation2:a
	signal memory_delay7_output_wire                                            : std_logic_vector(23 downto 0); -- Memory_Delay7:output -> cast112:input
	signal cast112_output_wire                                                  : std_logic_vector(40 downto 0); -- cast112:output -> Comparator:dataa
	signal comparator_result_wire                                               : std_logic;                     -- Comparator:result -> cast113:input
	signal cast113_output_wire                                                  : std_logic_vector(0 downto 0);  -- cast113:output -> Multiplexer:sel
	signal bus_conversion4_output_wire                                          : std_logic_vector(7 downto 0);  -- Bus_Conversion4:output -> cast114:input
	signal cast114_output_wire                                                  : std_logic_vector(15 downto 0); -- cast114:output -> Multiplexer:in0
	signal cast115_output_wire                                                  : std_logic_vector(7 downto 0);  -- cast115:output -> Multiplier:datab
	signal cast116_output_wire                                                  : std_logic_vector(39 downto 0); -- cast116:output -> Pipelined_Adder:dataa
	signal multiplier1_result_wire                                              : std_logic_vector(34 downto 0); -- Multiplier1:result -> cast117:input
	signal cast117_output_wire                                                  : std_logic_vector(39 downto 0); -- cast117:output -> Pipelined_Adder:datab
	signal clock_0_clock_output_clk                                             : std_logic;                     -- Clock_0:clock_out -> [Bus_Concatenation2:clock, Bus_Concatenation3:clock, Comparator:clock, Divider:clk, Memory_Delay1:clock, Memory_Delay2:clock, Memory_Delay3:clock, Memory_Delay4:clock, Memory_Delay5:clock, Memory_Delay6:clock, Memory_Delay7:clock, Memory_Delay9:clock, Multiplexer:clock, Multiplier1:clock, Multiplier:clock, Pipelined_Adder1:clock, Pipelined_Adder:clock, localedgepreserve_Fusion_Cal_A_B_2_Cal_MeanG_0:Clock, localedgepreserve_Fusion_Cal_A_B_2_Cal_MeanI_VarI_0:Clock, localedgepreserve_Fusion_Cal_A_B_2_generate_signals_0:Clock]
	signal clock_0_clock_output_reset                                           : std_logic;                     -- Clock_0:aclr_out -> [Bus_Concatenation2:aclr, Bus_Concatenation3:aclr, Comparator:sclr, Memory_Delay1:aclr, Memory_Delay2:aclr, Memory_Delay3:aclr, Memory_Delay4:aclr, Memory_Delay5:aclr, Memory_Delay6:aclr, Memory_Delay7:aclr, Memory_Delay9:aclr, Multiplexer:aclr, Multiplier1:aclr, Multiplier:aclr, Pipelined_Adder1:aclr, Pipelined_Adder:aclr, localedgepreserve_Fusion_Cal_A_B_2_Cal_MeanG_0:reset, localedgepreserve_Fusion_Cal_A_B_2_Cal_MeanI_VarI_0:reset, localedgepreserve_Fusion_Cal_A_B_2_generate_signals_0:reset]

begin

	clock_0 : component alt_dspbuilder_clock_GNQFU4PUDH
		port map (
			clock_out => clock_0_clock_output_clk,   -- clock_output.clk
			aclr_out  => clock_0_clock_output_reset, --             .reset
			clock     => Clock,                      --        clock.clk
			aclr      => reset                       --             .reset
		);

	valid_in_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => valid_in,               --  input.wire
			output => valid_in_0_output_wire  -- output.wire
		);

	multiplier1 : component alt_dspbuilder_multiplier_GN2GJCFTFE
		generic map (
			aWidth                         => 35,
			Signed                         => 0,
			bWidth                         => 24,
			DEDICATED_MULTIPLIER_CIRCUITRY => "YES",
			pipeline                       => 1,
			OutputLsb                      => 24,
			OutputMsb                      => 58
		)
		port map (
			clock     => clock_0_clock_output_clk,            -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,          --           .reset
			dataa     => memory_delay9_output_wire,           --      dataa.wire
			datab     => constant_1_output_wire,              --      datab.wire
			result    => multiplier1_result_wire,             --     result.wire
			user_aclr => multiplier1user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => valid_in_0_output_wire               --        ena.wire
		);

	multiplier1user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplier1user_aclrgnd_output_wire  -- output.wire
		);

	binary_point_casting1 : component alt_dspbuilder_cast_GNUYRTQ4QH
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => cast109_output_wire,               --  input.wire
			output => binary_point_casting1_output_wire  -- output.wire
		);

	eof_out_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => localedgepreserve_fusion_cal_a_b_2_generate_signals_0_eof_out_wire, --  input.wire
			output => eof_out                                                             -- output.wire
		);

	binary_point_casting3 : component alt_dspbuilder_cast_GNUYRTQ4QH
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => bus_conversion2_output_wire,       --  input.wire
			output => binary_point_casting3_output_wire  -- output.wire
		);

	binary_point_casting2 : component alt_dspbuilder_cast_GNUYRTQ4QH
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => bus_conversion3_output_wire,       --  input.wire
			output => binary_point_casting2_output_wire  -- output.wire
		);

	multiplexer : component alt_dspbuilder_multiplexer_GN7X7SG76C
		generic map (
			number_inputs          => 2,
			pipeline               => 0,
			width                  => 16,
			HDLTYPE                => "STD_LOGIC_VECTOR",
			use_one_hot_select_bus => 0
		)
		port map (
			clock     => clock_0_clock_output_clk,            -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,          --           .reset
			sel       => cast113_output_wire,                 --        sel.wire
			result    => multiplexer_result_wire,             --     result.wire
			ena       => multiplexerenavcc_output_wire,       --        ena.wire
			user_aclr => multiplexeruser_aclrgnd_output_wire, --  user_aclr.wire
			in0       => cast114_output_wire,                 --        in0.wire
			in1       => constant4_output_wire                --        in1.wire
		);

	multiplexeruser_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplexeruser_aclrgnd_output_wire  -- output.wire
		);

	multiplexerenavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => multiplexerenavcc_output_wire  -- output.wire
		);

	grad_in_0 : component alt_dspbuilder_port_GNLA26EJAH
		port map (
			input  => grad_in,               --  input.wire
			output => grad_in_0_output_wire  -- output.wire
		);

	pixel_in_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => pixel_in,               --  input.wire
			output => pixel_in_0_output_wire  -- output.wire
		);

	memory_delay7 : component alt_dspbuilder_memdelay_GNDI52L3LZ
		generic map (
			RAMTYPE => "AUTO",
			WIDTH   => 24,
			DELAY   => 25
		)
		port map (
			clock     => clock_0_clock_output_clk,              -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,            --           .reset
			input     => memory_delay2_output_wire,             --      input.wire
			output    => memory_delay7_output_wire,             --     output.wire
			user_aclr => memory_delay7user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => valid_in_0_output_wire                 --        ena.wire
		);

	memory_delay7user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => memory_delay7user_aclrgnd_output_wire  -- output.wire
		);

	pipelined_adder : component alt_dspbuilder_pipelined_adder_GNTWZRTG4I
		generic map (
			pipeline => 1,
			width    => 40
		)
		port map (
			clock     => clock_0_clock_output_clk,                -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,              --           .reset
			dataa     => cast116_output_wire,                     --      dataa.wire
			datab     => cast117_output_wire,                     --      datab.wire
			result    => pipelined_adder_result_wire,             --     result.wire
			user_aclr => pipelined_adderuser_aclrgnd_output_wire, --  user_aclr.wire
			ena       => valid_in_0_output_wire                   --        ena.wire
		);

	pipelined_adderuser_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => pipelined_adderuser_aclrgnd_output_wire  -- output.wire
		);

	memory_delay5 : component alt_dspbuilder_memdelay_GNMIZKWFE6
		generic map (
			RAMTYPE => "AUTO",
			WIDTH   => 16,
			DELAY   => 1
		)
		port map (
			clock     => clock_0_clock_output_clk,              -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,            --           .reset
			input     => memory_delay3_output_wire,             --      input.wire
			output    => memory_delay5_output_wire,             --     output.wire
			user_aclr => memory_delay5user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => valid_in_0_output_wire                 --        ena.wire
		);

	memory_delay5user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => memory_delay5user_aclrgnd_output_wire  -- output.wire
		);

	memory_delay6 : component alt_dspbuilder_memdelay_GNI6WYI4F7
		generic map (
			RAMTYPE => "AUTO",
			WIDTH   => 8,
			DELAY   => 29
		)
		port map (
			clock     => clock_0_clock_output_clk,                                           -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,                                         --           .reset
			input     => localedgepreserve_fusion_cal_a_b_2_cal_meani_vari_0_pixel_out_wire, --      input.wire
			output    => memory_delay6_output_wire,                                          --     output.wire
			user_aclr => memory_delay6user_aclrgnd_output_wire,                              --  user_aclr.wire
			ena       => valid_in_0_output_wire                                              --        ena.wire
		);

	memory_delay6user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => memory_delay6user_aclrgnd_output_wire  -- output.wire
		);

	localedgepreserve_fusion_cal_a_b_2_cal_meani_vari_0 : component localedgepreserve_GN_localedgepreserve_Fusion_Cal_A_B_2_Cal_MeanI_VarI
		port map (
			valid_in  => valid_in_0_output_wire,                                             --  valid_in.wire
			Clock     => clock_0_clock_output_clk,                                           --     Clock.clk
			reset     => clock_0_clock_output_reset,                                         --          .reset
			pixel_out => localedgepreserve_fusion_cal_a_b_2_cal_meani_vari_0_pixel_out_wire, -- pixel_out.wire
			pixel_in  => pixel_in_0_output_wire,                                             --  pixel_in.wire
			varI      => localedgepreserve_fusion_cal_a_b_2_cal_meani_vari_0_vari_wire,      --      varI.wire
			meanI     => localedgepreserve_fusion_cal_a_b_2_cal_meani_vari_0_meani_wire      --     meanI.wire
		);

	memory_delay9 : component alt_dspbuilder_memdelay_GNF7HJJOOI
		generic map (
			RAMTYPE => "AUTO",
			WIDTH   => 35,
			DELAY   => 2
		)
		port map (
			clock     => clock_0_clock_output_clk,                                  -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,                                --           .reset
			input     => localedgepreserve_fusion_cal_a_b_2_cal_meang_0_meang_wire, --      input.wire
			output    => memory_delay9_output_wire,                                 --     output.wire
			user_aclr => memory_delay9user_aclrgnd_output_wire,                     --  user_aclr.wire
			ena       => valid_in_0_output_wire                                     --        ena.wire
		);

	memory_delay9user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => memory_delay9user_aclrgnd_output_wire  -- output.wire
		);

	comparator : component alt_dspbuilder_comparator_GN
		generic map (
			Operator  => "Altaeb",
			lpm_width => 41
		)
		port map (
			clock  => clock_0_clock_output_clk,   -- clock_sclr.clk
			sclr   => clock_0_clock_output_reset, --           .reset
			dataa  => cast112_output_wire,        --      dataa.wire
			datab  => cast106_output_wire,        --      datab.wire
			result => comparator_result_wire      --     result.wire
		);

	valid_out_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => localedgepreserve_fusion_cal_a_b_2_generate_signals_0_valid_out_wire, --  input.wire
			output => valid_out                                                             -- output.wire
		);

	memory_delay3 : component alt_dspbuilder_memdelay_GN4TPDAUQN
		generic map (
			RAMTYPE => "AUTO",
			WIDTH   => 16,
			DELAY   => 27
		)
		port map (
			clock     => clock_0_clock_output_clk,              -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,            --           .reset
			input     => bus_conversion5_output_wire,           --      input.wire
			output    => memory_delay3_output_wire,             --     output.wire
			user_aclr => memory_delay3user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => valid_in_0_output_wire                 --        ena.wire
		);

	memory_delay3user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => memory_delay3user_aclrgnd_output_wire  -- output.wire
		);

	memory_delay4 : component alt_dspbuilder_memdelay_GNMYXI7BAD
		generic map (
			RAMTYPE => "AUTO",
			WIDTH   => 16,
			DELAY   => 2
		)
		port map (
			clock     => clock_0_clock_output_clk,              -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,            --           .reset
			input     => multiplexer_result_wire,               --      input.wire
			output    => memory_delay4_output_wire,             --     output.wire
			user_aclr => memory_delay4user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => valid_in_0_output_wire                 --        ena.wire
		);

	memory_delay4user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => memory_delay4user_aclrgnd_output_wire  -- output.wire
		);

	memory_delay1 : component alt_dspbuilder_memdelay_GNNY7HWC5A
		generic map (
			RAMTYPE => "AUTO",
			WIDTH   => 40,
			DELAY   => 1
		)
		port map (
			clock     => clock_0_clock_output_clk,                                      -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,                                    --           .reset
			input     => localedgepreserve_fusion_cal_a_b_2_cal_meani_vari_0_vari_wire, --      input.wire
			output    => memory_delay1_output_wire,                                     --     output.wire
			user_aclr => memory_delay1user_aclrgnd_output_wire,                         --  user_aclr.wire
			ena       => valid_in_0_output_wire                                         --        ena.wire
		);

	memory_delay1user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => memory_delay1user_aclrgnd_output_wire  -- output.wire
		);

	memory_delay2 : component alt_dspbuilder_memdelay_GNZWVQQT43
		generic map (
			RAMTYPE => "AUTO",
			WIDTH   => 24,
			DELAY   => 1
		)
		port map (
			clock     => clock_0_clock_output_clk,              -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,            --           .reset
			input     => binary_point_casting3_output_wire,     --      input.wire
			output    => memory_delay2_output_wire,             --     output.wire
			user_aclr => memory_delay2user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => valid_in_0_output_wire                 --        ena.wire
		);

	memory_delay2user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => memory_delay2user_aclrgnd_output_wire  -- output.wire
		);

	multiplier : component alt_dspbuilder_multiplier_GNKTEWW72G
		generic map (
			aWidth                         => 16,
			Signed                         => 0,
			bWidth                         => 8,
			DEDICATED_MULTIPLIER_CIRCUITRY => "YES",
			pipeline                       => 1,
			OutputLsb                      => 8,
			OutputMsb                      => 23
		)
		port map (
			clock     => clock_0_clock_output_clk,           -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,         --           .reset
			dataa     => memory_delay3_output_wire,          --      dataa.wire
			datab     => cast115_output_wire,                --      datab.wire
			result    => multiplier_result_wire,             --     result.wire
			user_aclr => multiplieruser_aclrgnd_output_wire, --  user_aclr.wire
			ena       => valid_in_0_output_wire              --        ena.wire
		);

	multiplieruser_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplieruser_aclrgnd_output_wire  -- output.wire
		);

	pipelined_adder1 : component alt_dspbuilder_pipelined_adder_GNWEIMU3MK
		generic map (
			pipeline => 1,
			width    => 16
		)
		port map (
			clock     => clock_0_clock_output_clk,                 -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,               --           .reset
			dataa     => memory_delay5_output_wire,                --      dataa.wire
			datab     => multiplier_result_wire,                   --      datab.wire
			result    => pipelined_adder1_result_wire,             --     result.wire
			user_aclr => pipelined_adder1user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => valid_in_0_output_wire                    --        ena.wire
		);

	pipelined_adder1user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => pipelined_adder1user_aclrgnd_output_wire  -- output.wire
		);

	bus_conversion5 : component alt_dspbuilder_cast_GNPPZDVXTY
		generic map (
			round    => 1,
			saturate => 0
		)
		port map (
			input  => localedgepreserve_fusion_cal_a_b_2_cal_meani_vari_0_meani_wire, --  input.wire
			output => bus_conversion5_output_wire                                     -- output.wire
		);

	bus_conversion4 : component alt_dspbuilder_cast_GNW6I55EUT
		generic map (
			round    => 1,
			saturate => 0
		)
		port map (
			input  => binary_point_casting1_output_wire, --  input.wire
			output => bus_conversion4_output_wire        -- output.wire
		);

	b_out_0 : component alt_dspbuilder_port_GNBO6OMO5Y
		port map (
			input  => pipelined_adder1_result_wire, --  input.wire
			output => b_out                         -- output.wire
		);

	bus_conversion3 : component alt_dspbuilder_cast_GNZYD62DLY
		generic map (
			round    => 1,
			saturate => 0
		)
		port map (
			input  => pipelined_adder_result_wire, --  input.wire
			output => bus_conversion3_output_wire  -- output.wire
		);

	bus_conversion2 : component alt_dspbuilder_cast_GNZYD62DLY
		generic map (
			round    => 1,
			saturate => 0
		)
		port map (
			input  => cast110_output_wire,         --  input.wire
			output => bus_conversion2_output_wire  -- output.wire
		);

	localedgepreserve_fusion_cal_a_b_2_cal_meang_0 : component localedgepreserve_GN_localedgepreserve_Fusion_Cal_A_B_2_Cal_MeanG
		port map (
			meanG    => localedgepreserve_fusion_cal_a_b_2_cal_meang_0_meang_wire, --    meanG.wire
			Clock    => clock_0_clock_output_clk,                                  --    Clock.clk
			reset    => clock_0_clock_output_reset,                                --         .reset
			valid_in => valid_in_0_output_wire,                                    -- valid_in.wire
			pixel_in => grad_in_0_output_wire                                      -- pixel_in.wire
		);

	constant1 : component alt_dspbuilder_constant_GNRSDUIWRP
		generic map (
			BitPattern => "00000000000000000000000000000000",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 32
		)
		port map (
			output => constant1_output_wire  -- output.wire
		);

	localedgepreserve_fusion_cal_a_b_2_generate_signals_0 : component localedgepreserve_GN_localedgepreserve_Fusion_Cal_A_B_2_generate_signals
		port map (
			Clock     => clock_0_clock_output_clk,                                             --     Clock.clk
			reset     => clock_0_clock_output_reset,                                           --          .reset
			valid_in  => valid_in_0_output_wire,                                               --  valid_in.wire
			eof_out   => localedgepreserve_fusion_cal_a_b_2_generate_signals_0_eof_out_wire,   --   eof_out.wire
			valid_out => localedgepreserve_fusion_cal_a_b_2_generate_signals_0_valid_out_wire, -- valid_out.wire
			eof_in    => eof_in_0_output_wire                                                  --    eof_in.wire
		);

	eof_in_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => eof_in,               --  input.wire
			output => eof_in_0_output_wire  -- output.wire
		);

	bus_concatenation2 : component alt_dspbuilder_bus_concat_GNOQTN4QAD
		generic map (
			widthA => 24,
			widthB => 8
		)
		port map (
			clock  => clock_0_clock_output_clk,       -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,     --           .reset
			a      => cast111_output_wire,            --          a.wire
			b      => constant6_output_wire,          --          b.wire
			output => bus_concatenation2_output_wire  --     output.wire
		);

	bus_concatenation3 : component alt_dspbuilder_bus_concat_GNDDREGCTK
		generic map (
			widthA => 16,
			widthB => 32
		)
		port map (
			clock  => clock_0_clock_output_clk,       -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,     --           .reset
			a      => constant7_output_wire,          --          a.wire
			b      => bus_concatenation2_output_wire, --          b.wire
			output => bus_concatenation3_output_wire  --     output.wire
		);

	a_out_0 : component alt_dspbuilder_port_GNBO6OMO5Y
		port map (
			input  => memory_delay4_output_wire, --  input.wire
			output => a_out                      -- output.wire
		);

	constant6 : component alt_dspbuilder_constant_GNC5NOVIJT
		generic map (
			BitPattern => "00000000",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 8
		)
		port map (
			output => constant6_output_wire  -- output.wire
		);

	constant7 : component alt_dspbuilder_constant_GNCWI5QDAD
		generic map (
			BitPattern => "0000000000000000",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 16
		)
		port map (
			output => constant7_output_wire  -- output.wire
		);

	constant4 : component alt_dspbuilder_constant_GNCWI5QDAD
		generic map (
			BitPattern => "0000000000000000",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 16
		)
		port map (
			output => constant4_output_wire  -- output.wire
		);

	constant_1 : component alt_dspbuilder_constant_GN5FET4EJH
		generic map (
			BitPattern => "000110011001100110011001",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 24
		)
		port map (
			output => constant_1_output_wire  -- output.wire
		);

	pixel_out_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => memory_delay6_output_wire, --  input.wire
			output => pixel_out                  -- output.wire
		);

	divider : component div
		port map (
			clk => clock_0_clock_output_clk, -- clk.clk
			ena => valid_in_0_output_wire,   -- ena.wire
			z   => cast107_output_wire,      --   z.wire
			d   => cast108_output_wire,      --   d.wire
			q   => divider_q_wire            --   q.wire
		);

	cast106 : component alt_dspbuilder_cast_GN3FODBL3U
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => constant1_output_wire, --  input.wire
			output => cast106_output_wire    -- output.wire
		);

	cast107 : component alt_dspbuilder_cast_GNKD3JEUSD
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => bus_concatenation3_output_wire, --  input.wire
			output => cast107_output_wire             -- output.wire
		);

	cast108 : component alt_dspbuilder_cast_GN5P6ORZXA
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => binary_point_casting2_output_wire, --  input.wire
			output => cast108_output_wire                -- output.wire
		);

	cast109 : component alt_dspbuilder_cast_GNEIIG67TZ
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => divider_q_wire,      --  input.wire
			output => cast109_output_wire  -- output.wire
		);

	cast110 : component alt_dspbuilder_cast_GNOEMJJSIT
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => memory_delay1_output_wire, --  input.wire
			output => cast110_output_wire        -- output.wire
		);

	cast111 : component alt_dspbuilder_cast_GNA5TAMWCZ
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => memory_delay2_output_wire, --  input.wire
			output => cast111_output_wire        -- output.wire
		);

	cast112 : component alt_dspbuilder_cast_GNP5J2CFQQ
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => memory_delay7_output_wire, --  input.wire
			output => cast112_output_wire        -- output.wire
		);

	cast113 : component alt_dspbuilder_cast_GN46N4UJ5S
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => comparator_result_wire, --  input.wire
			output => cast113_output_wire     -- output.wire
		);

	cast114 : component alt_dspbuilder_cast_GNDHESB5KA
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => bus_conversion4_output_wire, --  input.wire
			output => cast114_output_wire          -- output.wire
		);

	cast115 : component alt_dspbuilder_cast_GNT7Y2ULVV
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => multiplexer_result_wire, --  input.wire
			output => cast115_output_wire      -- output.wire
		);

	cast116 : component alt_dspbuilder_cast_GNOEMJJSIT
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => memory_delay1_output_wire, --  input.wire
			output => cast116_output_wire        -- output.wire
		);

	cast117 : component alt_dspbuilder_cast_GNXSA7APAK
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => multiplier1_result_wire, --  input.wire
			output => cast117_output_wire      -- output.wire
		);

end architecture rtl; -- of localedgepreserve_GN_localedgepreserve_Fusion_Cal_A_B_2
