// de2i_150_qsys.v

// Generated using ACDS version 17.1 590

`timescale 1 ps / 1 ps
module de2i_150_qsys (
		input  wire        alt_vip_itc_0_clocked_video_vid_clk,        // alt_vip_itc_0_clocked_video.vid_clk
		output wire [23:0] alt_vip_itc_0_clocked_video_vid_data,       //                            .vid_data
		output wire        alt_vip_itc_0_clocked_video_underflow,      //                            .underflow
		output wire        alt_vip_itc_0_clocked_video_vid_datavalid,  //                            .vid_datavalid
		output wire        alt_vip_itc_0_clocked_video_vid_v_sync,     //                            .vid_v_sync
		output wire        alt_vip_itc_0_clocked_video_vid_h_sync,     //                            .vid_h_sync
		output wire        alt_vip_itc_0_clocked_video_vid_f,          //                            .vid_f
		output wire        alt_vip_itc_0_clocked_video_vid_h,          //                            .vid_h
		output wire        alt_vip_itc_0_clocked_video_vid_v,          //                            .vid_v
		output wire        altpll_sdram_clk,                           //                altpll_sdram.clk
		output wire        altpll_vga_clk,                             //                  altpll_vga.clk
		input  wire        clk_clk,                                    //                         clk.clk
		output wire        pcie_ip_clocks_sim_clk250_export,           //          pcie_ip_clocks_sim.clk250_export
		output wire        pcie_ip_clocks_sim_clk500_export,           //                            .clk500_export
		output wire        pcie_ip_clocks_sim_clk125_export,           //                            .clk125_export
		input  wire        pcie_ip_pcie_rstn_export,                   //           pcie_ip_pcie_rstn.export
		input  wire        pcie_ip_pipe_ext_pipe_mode,                 //            pcie_ip_pipe_ext.pipe_mode
		input  wire        pcie_ip_pipe_ext_phystatus_ext,             //                            .phystatus_ext
		output wire        pcie_ip_pipe_ext_rate_ext,                  //                            .rate_ext
		output wire [1:0]  pcie_ip_pipe_ext_powerdown_ext,             //                            .powerdown_ext
		output wire        pcie_ip_pipe_ext_txdetectrx_ext,            //                            .txdetectrx_ext
		input  wire        pcie_ip_pipe_ext_rxelecidle0_ext,           //                            .rxelecidle0_ext
		input  wire [7:0]  pcie_ip_pipe_ext_rxdata0_ext,               //                            .rxdata0_ext
		input  wire [2:0]  pcie_ip_pipe_ext_rxstatus0_ext,             //                            .rxstatus0_ext
		input  wire        pcie_ip_pipe_ext_rxvalid0_ext,              //                            .rxvalid0_ext
		input  wire        pcie_ip_pipe_ext_rxdatak0_ext,              //                            .rxdatak0_ext
		output wire [7:0]  pcie_ip_pipe_ext_txdata0_ext,               //                            .txdata0_ext
		output wire        pcie_ip_pipe_ext_txdatak0_ext,              //                            .txdatak0_ext
		output wire        pcie_ip_pipe_ext_rxpolarity0_ext,           //                            .rxpolarity0_ext
		output wire        pcie_ip_pipe_ext_txcompl0_ext,              //                            .txcompl0_ext
		output wire        pcie_ip_pipe_ext_txelecidle0_ext,           //                            .txelecidle0_ext
		input  wire        pcie_ip_reconfig_busy_busy_altgxb_reconfig, //       pcie_ip_reconfig_busy.busy_altgxb_reconfig
		output wire [4:0]  pcie_ip_reconfig_fromgxb_0_data,            //  pcie_ip_reconfig_fromgxb_0.data
		input  wire [3:0]  pcie_ip_reconfig_togxb_data,                //      pcie_ip_reconfig_togxb.data
		input  wire        pcie_ip_refclk_export,                      //              pcie_ip_refclk.export
		input  wire        pcie_ip_rx_in_rx_datain_0,                  //               pcie_ip_rx_in.rx_datain_0
		input  wire [39:0] pcie_ip_test_in_test_in,                    //             pcie_ip_test_in.test_in
		output wire        pcie_ip_tx_out_tx_dataout_0,                //              pcie_ip_tx_out.tx_dataout_0
		input  wire        reset_reset_n,                              //                       reset.reset_n
		output wire [12:0] sdram_addr,                                 //                       sdram.addr
		output wire [1:0]  sdram_ba,                                   //                            .ba
		output wire        sdram_cas_n,                                //                            .cas_n
		output wire        sdram_cke,                                  //                            .cke
		output wire        sdram_cs_n,                                 //                            .cs_n
		inout  wire [31:0] sdram_dq,                                   //                            .dq
		output wire [3:0]  sdram_dqm,                                  //                            .dqm
		output wire        sdram_ras_n,                                //                            .ras_n
		output wire        sdram_we_n,                                 //                            .we_n
		input  wire [1:0]  switch_name                                 //                      switch.name
	);

	wire          dma_read_master_data_source_valid;                                       // dma_read_master:src_valid -> dma_write_master:snk_valid
	wire   [31:0] dma_read_master_data_source_data;                                        // dma_read_master:src_data -> dma_write_master:snk_data
	wire          dma_read_master_data_source_ready;                                       // dma_write_master:snk_ready -> dma_read_master:src_ready
	wire          modular_sgdma_dispatcher_read_command_source_valid;                      // modular_sgdma_dispatcher:src_read_master_valid -> dma_read_master:snk_command_valid
	wire  [255:0] modular_sgdma_dispatcher_read_command_source_data;                       // modular_sgdma_dispatcher:src_read_master_data -> dma_read_master:snk_command_data
	wire          modular_sgdma_dispatcher_read_command_source_ready;                      // dma_read_master:snk_command_ready -> modular_sgdma_dispatcher:src_read_master_ready
	wire          dma_read_master_response_source_valid;                                   // dma_read_master:src_response_valid -> modular_sgdma_dispatcher:snk_read_master_valid
	wire  [255:0] dma_read_master_response_source_data;                                    // dma_read_master:src_response_data -> modular_sgdma_dispatcher:snk_read_master_data
	wire          dma_read_master_response_source_ready;                                   // modular_sgdma_dispatcher:snk_read_master_ready -> dma_read_master:src_response_ready
	wire          dma_write_master_response_source_valid;                                  // dma_write_master:src_response_valid -> modular_sgdma_dispatcher:snk_write_master_valid
	wire  [255:0] dma_write_master_response_source_data;                                   // dma_write_master:src_response_data -> modular_sgdma_dispatcher:snk_write_master_data
	wire          dma_write_master_response_source_ready;                                  // modular_sgdma_dispatcher:snk_write_master_ready -> dma_write_master:src_response_ready
	wire          modular_sgdma_dispatcher_write_command_source_valid;                     // modular_sgdma_dispatcher:src_write_master_valid -> dma_write_master:snk_command_valid
	wire  [255:0] modular_sgdma_dispatcher_write_command_source_data;                      // modular_sgdma_dispatcher:src_write_master_data -> dma_write_master:snk_command_data
	wire          modular_sgdma_dispatcher_write_command_source_ready;                     // dma_write_master:snk_command_ready -> modular_sgdma_dispatcher:src_write_master_ready
	wire          image1_padding_avalon_clipper_source_valid;                              // image1_padding:stream_out_valid -> image_fusion:sink1_valid
	wire    [7:0] image1_padding_avalon_clipper_source_data;                               // image1_padding:stream_out_data -> image_fusion:sink1_data
	wire          image1_padding_avalon_clipper_source_ready;                              // image_fusion:sink1_ready -> image1_padding:stream_out_ready
	wire          image1_padding_avalon_clipper_source_startofpacket;                      // image1_padding:stream_out_startofpacket -> image_fusion:sink1_sop
	wire          image1_padding_avalon_clipper_source_endofpacket;                        // image1_padding:stream_out_endofpacket -> image_fusion:sink1_eop
	wire          image2_padding_avalon_clipper_source_valid;                              // image2_padding:stream_out_valid -> image_fusion:sink2_valid
	wire    [7:0] image2_padding_avalon_clipper_source_data;                               // image2_padding:stream_out_data -> image_fusion:sink2_data
	wire          image2_padding_avalon_clipper_source_ready;                              // image_fusion:sink2_ready -> image2_padding:stream_out_ready
	wire          image2_padding_avalon_clipper_source_startofpacket;                      // image2_padding:stream_out_startofpacket -> image_fusion:sink2_sop
	wire          image2_padding_avalon_clipper_source_endofpacket;                        // image2_padding:stream_out_endofpacket -> image_fusion:sink2_eop
	wire          video_dma1_read_avalon_pixel_source_valid;                               // video_dma1_read:stream_valid -> buffer1_read:in_valid
	wire    [7:0] video_dma1_read_avalon_pixel_source_data;                                // video_dma1_read:stream_data -> buffer1_read:in_data
	wire          video_dma1_read_avalon_pixel_source_ready;                               // buffer1_read:in_ready -> video_dma1_read:stream_ready
	wire          video_dma1_read_avalon_pixel_source_startofpacket;                       // video_dma1_read:stream_startofpacket -> buffer1_read:in_startofpacket
	wire          video_dma1_read_avalon_pixel_source_endofpacket;                         // video_dma1_read:stream_endofpacket -> buffer1_read:in_endofpacket
	wire          video_dma2_read_avalon_pixel_source_valid;                               // video_dma2_read:stream_valid -> buffer2_read:in_valid
	wire    [7:0] video_dma2_read_avalon_pixel_source_data;                                // video_dma2_read:stream_data -> buffer2_read:in_data
	wire          video_dma2_read_avalon_pixel_source_ready;                               // buffer2_read:in_ready -> video_dma2_read:stream_ready
	wire          video_dma2_read_avalon_pixel_source_startofpacket;                       // video_dma2_read:stream_startofpacket -> buffer2_read:in_startofpacket
	wire          video_dma2_read_avalon_pixel_source_endofpacket;                         // video_dma2_read:stream_endofpacket -> buffer2_read:in_endofpacket
	wire          alt_vip_vfr_0_avalon_streaming_source_valid;                             // alt_vip_vfr_0:dout_valid -> alt_vip_itc_0:is_valid
	wire   [23:0] alt_vip_vfr_0_avalon_streaming_source_data;                              // alt_vip_vfr_0:dout_data -> alt_vip_itc_0:is_data
	wire          alt_vip_vfr_0_avalon_streaming_source_ready;                             // alt_vip_itc_0:is_ready -> alt_vip_vfr_0:dout_ready
	wire          alt_vip_vfr_0_avalon_streaming_source_startofpacket;                     // alt_vip_vfr_0:dout_startofpacket -> alt_vip_itc_0:is_sop
	wire          alt_vip_vfr_0_avalon_streaming_source_endofpacket;                       // alt_vip_vfr_0:dout_endofpacket -> alt_vip_itc_0:is_eop
	wire          buffer1_read_out_valid;                                                  // buffer1_read:out_valid -> image1_padding:stream_in_valid
	wire    [7:0] buffer1_read_out_data;                                                   // buffer1_read:out_data -> image1_padding:stream_in_data
	wire          buffer1_read_out_ready;                                                  // image1_padding:stream_in_ready -> buffer1_read:out_ready
	wire          buffer1_read_out_startofpacket;                                          // buffer1_read:out_startofpacket -> image1_padding:stream_in_startofpacket
	wire          buffer1_read_out_endofpacket;                                            // buffer1_read:out_endofpacket -> image1_padding:stream_in_endofpacket
	wire          buffer2_read_out_valid;                                                  // buffer2_read:out_valid -> image2_padding:stream_in_valid
	wire    [7:0] buffer2_read_out_data;                                                   // buffer2_read:out_data -> image2_padding:stream_in_data
	wire          buffer2_read_out_ready;                                                  // image2_padding:stream_in_ready -> buffer2_read:out_ready
	wire          buffer2_read_out_startofpacket;                                          // buffer2_read:out_startofpacket -> image2_padding:stream_in_startofpacket
	wire          buffer2_read_out_endofpacket;                                            // buffer2_read:out_endofpacket -> image2_padding:stream_in_endofpacket
	wire          altpll_qsys_c0_clk;                                                      // altpll_qsys:c0 -> [alt_vip_itc_0:is_clk, alt_vip_vfr_0:clock, alt_vip_vfr_0:master_clock, avalon_st_adapter:in_clk_0_clk, avalon_st_adapter_001:in_clk_0_clk, buffer1_read:clk, buffer2_read:clk, buffer_write:clk, image1_padding:clk, image2_padding:clk, image_fusion:Clock, mm_interconnect_0:altpll_qsys_c0_clk, mm_interconnect_1:altpll_qsys_c0_clk, rst_controller:clk, sdram:clk, video_dma1_read:clk, video_dma2_read:clk, video_dma_write:clk]
	wire          altpll_qsys_c3_clk;                                                      // altpll_qsys:c3 -> [pcie_ip:cal_blk_clk_clk, pcie_ip:reconfig_gxbclk_clk]
	wire          pcie_ip_pcie_core_clk_clk;                                               // pcie_ip:pcie_core_clk_clk -> [dma_read_master:clk, dma_write_master:clk, irq_mapper:clk, mm_interconnect_0:pcie_ip_pcie_core_clk_clk, mm_interconnect_1:pcie_ip_pcie_core_clk_clk, mm_interconnect_2:pcie_ip_pcie_core_clk_clk, modular_sgdma_dispatcher:clk, pcie_ip:fixedclk_clk, rst_controller_002:clk]
	wire   [31:0] dma_read_master_data_read_master_readdata;                               // mm_interconnect_0:dma_read_master_Data_Read_Master_readdata -> dma_read_master:master_readdata
	wire          dma_read_master_data_read_master_waitrequest;                            // mm_interconnect_0:dma_read_master_Data_Read_Master_waitrequest -> dma_read_master:master_waitrequest
	wire   [31:0] dma_read_master_data_read_master_address;                                // dma_read_master:master_address -> mm_interconnect_0:dma_read_master_Data_Read_Master_address
	wire          dma_read_master_data_read_master_read;                                   // dma_read_master:master_read -> mm_interconnect_0:dma_read_master_Data_Read_Master_read
	wire    [3:0] dma_read_master_data_read_master_byteenable;                             // dma_read_master:master_byteenable -> mm_interconnect_0:dma_read_master_Data_Read_Master_byteenable
	wire          dma_read_master_data_read_master_readdatavalid;                          // mm_interconnect_0:dma_read_master_Data_Read_Master_readdatavalid -> dma_read_master:master_readdatavalid
	wire    [4:0] dma_read_master_data_read_master_burstcount;                             // dma_read_master:master_burstcount -> mm_interconnect_0:dma_read_master_Data_Read_Master_burstcount
	wire          dma_write_master_data_write_master_waitrequest;                          // mm_interconnect_0:dma_write_master_Data_Write_Master_waitrequest -> dma_write_master:master_waitrequest
	wire   [31:0] dma_write_master_data_write_master_address;                              // dma_write_master:master_address -> mm_interconnect_0:dma_write_master_Data_Write_Master_address
	wire    [3:0] dma_write_master_data_write_master_byteenable;                           // dma_write_master:master_byteenable -> mm_interconnect_0:dma_write_master_Data_Write_Master_byteenable
	wire          dma_write_master_data_write_master_write;                                // dma_write_master:master_write -> mm_interconnect_0:dma_write_master_Data_Write_Master_write
	wire   [31:0] dma_write_master_data_write_master_writedata;                            // dma_write_master:master_writedata -> mm_interconnect_0:dma_write_master_Data_Write_Master_writedata
	wire    [4:0] dma_write_master_data_write_master_burstcount;                           // dma_write_master:master_burstcount -> mm_interconnect_0:dma_write_master_Data_Write_Master_burstcount
	wire          video_dma1_read_avalon_dma_master_waitrequest;                           // mm_interconnect_0:video_dma1_read_avalon_dma_master_waitrequest -> video_dma1_read:master_waitrequest
	wire    [7:0] video_dma1_read_avalon_dma_master_readdata;                              // mm_interconnect_0:video_dma1_read_avalon_dma_master_readdata -> video_dma1_read:master_readdata
	wire   [31:0] video_dma1_read_avalon_dma_master_address;                               // video_dma1_read:master_address -> mm_interconnect_0:video_dma1_read_avalon_dma_master_address
	wire          video_dma1_read_avalon_dma_master_read;                                  // video_dma1_read:master_read -> mm_interconnect_0:video_dma1_read_avalon_dma_master_read
	wire          video_dma1_read_avalon_dma_master_readdatavalid;                         // mm_interconnect_0:video_dma1_read_avalon_dma_master_readdatavalid -> video_dma1_read:master_readdatavalid
	wire          video_dma1_read_avalon_dma_master_lock;                                  // video_dma1_read:master_arbiterlock -> mm_interconnect_0:video_dma1_read_avalon_dma_master_lock
	wire          video_dma_write_avalon_dma_master_waitrequest;                           // mm_interconnect_0:video_dma_write_avalon_dma_master_waitrequest -> video_dma_write:master_waitrequest
	wire   [31:0] video_dma_write_avalon_dma_master_address;                               // video_dma_write:master_address -> mm_interconnect_0:video_dma_write_avalon_dma_master_address
	wire          video_dma_write_avalon_dma_master_write;                                 // video_dma_write:master_write -> mm_interconnect_0:video_dma_write_avalon_dma_master_write
	wire   [31:0] video_dma_write_avalon_dma_master_writedata;                             // video_dma_write:master_writedata -> mm_interconnect_0:video_dma_write_avalon_dma_master_writedata
	wire          video_dma2_read_avalon_dma_master_waitrequest;                           // mm_interconnect_0:video_dma2_read_avalon_dma_master_waitrequest -> video_dma2_read:master_waitrequest
	wire    [7:0] video_dma2_read_avalon_dma_master_readdata;                              // mm_interconnect_0:video_dma2_read_avalon_dma_master_readdata -> video_dma2_read:master_readdata
	wire   [31:0] video_dma2_read_avalon_dma_master_address;                               // video_dma2_read:master_address -> mm_interconnect_0:video_dma2_read_avalon_dma_master_address
	wire          video_dma2_read_avalon_dma_master_read;                                  // video_dma2_read:master_read -> mm_interconnect_0:video_dma2_read_avalon_dma_master_read
	wire          video_dma2_read_avalon_dma_master_readdatavalid;                         // mm_interconnect_0:video_dma2_read_avalon_dma_master_readdatavalid -> video_dma2_read:master_readdatavalid
	wire          video_dma2_read_avalon_dma_master_lock;                                  // video_dma2_read:master_arbiterlock -> mm_interconnect_0:video_dma2_read_avalon_dma_master_lock
	wire   [31:0] alt_vip_vfr_0_avalon_master_readdata;                                    // mm_interconnect_0:alt_vip_vfr_0_avalon_master_readdata -> alt_vip_vfr_0:master_readdata
	wire          alt_vip_vfr_0_avalon_master_waitrequest;                                 // mm_interconnect_0:alt_vip_vfr_0_avalon_master_waitrequest -> alt_vip_vfr_0:master_waitrequest
	wire   [31:0] alt_vip_vfr_0_avalon_master_address;                                     // alt_vip_vfr_0:master_address -> mm_interconnect_0:alt_vip_vfr_0_avalon_master_address
	wire          alt_vip_vfr_0_avalon_master_read;                                        // alt_vip_vfr_0:master_read -> mm_interconnect_0:alt_vip_vfr_0_avalon_master_read
	wire          alt_vip_vfr_0_avalon_master_readdatavalid;                               // mm_interconnect_0:alt_vip_vfr_0_avalon_master_readdatavalid -> alt_vip_vfr_0:master_readdatavalid
	wire    [5:0] alt_vip_vfr_0_avalon_master_burstcount;                                  // alt_vip_vfr_0:master_burstcount -> mm_interconnect_0:alt_vip_vfr_0_avalon_master_burstcount
	wire          mm_interconnect_0_sdram_s1_chipselect;                                   // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire   [31:0] mm_interconnect_0_sdram_s1_readdata;                                     // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire          mm_interconnect_0_sdram_s1_waitrequest;                                  // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire   [24:0] mm_interconnect_0_sdram_s1_address;                                      // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire          mm_interconnect_0_sdram_s1_read;                                         // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire    [3:0] mm_interconnect_0_sdram_s1_byteenable;                                   // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire          mm_interconnect_0_sdram_s1_readdatavalid;                                // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire          mm_interconnect_0_sdram_s1_write;                                        // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire   [31:0] mm_interconnect_0_sdram_s1_writedata;                                    // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire          mm_interconnect_0_pcie_ip_txs_chipselect;                                // mm_interconnect_0:pcie_ip_txs_chipselect -> pcie_ip:txs_chipselect
	wire   [63:0] mm_interconnect_0_pcie_ip_txs_readdata;                                  // pcie_ip:txs_readdata -> mm_interconnect_0:pcie_ip_txs_readdata
	wire          mm_interconnect_0_pcie_ip_txs_waitrequest;                               // pcie_ip:txs_waitrequest -> mm_interconnect_0:pcie_ip_txs_waitrequest
	wire   [30:0] mm_interconnect_0_pcie_ip_txs_address;                                   // mm_interconnect_0:pcie_ip_txs_address -> pcie_ip:txs_address
	wire          mm_interconnect_0_pcie_ip_txs_read;                                      // mm_interconnect_0:pcie_ip_txs_read -> pcie_ip:txs_read
	wire    [7:0] mm_interconnect_0_pcie_ip_txs_byteenable;                                // mm_interconnect_0:pcie_ip_txs_byteenable -> pcie_ip:txs_byteenable
	wire          mm_interconnect_0_pcie_ip_txs_readdatavalid;                             // pcie_ip:txs_readdatavalid -> mm_interconnect_0:pcie_ip_txs_readdatavalid
	wire          mm_interconnect_0_pcie_ip_txs_write;                                     // mm_interconnect_0:pcie_ip_txs_write -> pcie_ip:txs_write
	wire   [63:0] mm_interconnect_0_pcie_ip_txs_writedata;                                 // mm_interconnect_0:pcie_ip_txs_writedata -> pcie_ip:txs_writedata
	wire    [6:0] mm_interconnect_0_pcie_ip_txs_burstcount;                                // mm_interconnect_0:pcie_ip_txs_burstcount -> pcie_ip:txs_burstcount
	wire          pcie_ip_bar1_0_waitrequest;                                              // mm_interconnect_1:pcie_ip_bar1_0_waitrequest -> pcie_ip:bar1_0_waitrequest
	wire   [63:0] pcie_ip_bar1_0_readdata;                                                 // mm_interconnect_1:pcie_ip_bar1_0_readdata -> pcie_ip:bar1_0_readdata
	wire   [31:0] pcie_ip_bar1_0_address;                                                  // pcie_ip:bar1_0_address -> mm_interconnect_1:pcie_ip_bar1_0_address
	wire          pcie_ip_bar1_0_read;                                                     // pcie_ip:bar1_0_read -> mm_interconnect_1:pcie_ip_bar1_0_read
	wire    [7:0] pcie_ip_bar1_0_byteenable;                                               // pcie_ip:bar1_0_byteenable -> mm_interconnect_1:pcie_ip_bar1_0_byteenable
	wire          pcie_ip_bar1_0_readdatavalid;                                            // mm_interconnect_1:pcie_ip_bar1_0_readdatavalid -> pcie_ip:bar1_0_readdatavalid
	wire          pcie_ip_bar1_0_write;                                                    // pcie_ip:bar1_0_write -> mm_interconnect_1:pcie_ip_bar1_0_write
	wire   [63:0] pcie_ip_bar1_0_writedata;                                                // pcie_ip:bar1_0_writedata -> mm_interconnect_1:pcie_ip_bar1_0_writedata
	wire    [6:0] pcie_ip_bar1_0_burstcount;                                               // pcie_ip:bar1_0_burstcount -> mm_interconnect_1:pcie_ip_bar1_0_burstcount
	wire   [31:0] mm_interconnect_1_video_dma_write_avalon_dma_control_slave_readdata;     // video_dma_write:slave_readdata -> mm_interconnect_1:video_dma_write_avalon_dma_control_slave_readdata
	wire    [1:0] mm_interconnect_1_video_dma_write_avalon_dma_control_slave_address;      // mm_interconnect_1:video_dma_write_avalon_dma_control_slave_address -> video_dma_write:slave_address
	wire          mm_interconnect_1_video_dma_write_avalon_dma_control_slave_read;         // mm_interconnect_1:video_dma_write_avalon_dma_control_slave_read -> video_dma_write:slave_read
	wire    [3:0] mm_interconnect_1_video_dma_write_avalon_dma_control_slave_byteenable;   // mm_interconnect_1:video_dma_write_avalon_dma_control_slave_byteenable -> video_dma_write:slave_byteenable
	wire          mm_interconnect_1_video_dma_write_avalon_dma_control_slave_write;        // mm_interconnect_1:video_dma_write_avalon_dma_control_slave_write -> video_dma_write:slave_write
	wire   [31:0] mm_interconnect_1_video_dma_write_avalon_dma_control_slave_writedata;    // mm_interconnect_1:video_dma_write_avalon_dma_control_slave_writedata -> video_dma_write:slave_writedata
	wire   [31:0] mm_interconnect_1_video_dma1_read_avalon_dma_control_slave_readdata;     // video_dma1_read:slave_readdata -> mm_interconnect_1:video_dma1_read_avalon_dma_control_slave_readdata
	wire    [1:0] mm_interconnect_1_video_dma1_read_avalon_dma_control_slave_address;      // mm_interconnect_1:video_dma1_read_avalon_dma_control_slave_address -> video_dma1_read:slave_address
	wire          mm_interconnect_1_video_dma1_read_avalon_dma_control_slave_read;         // mm_interconnect_1:video_dma1_read_avalon_dma_control_slave_read -> video_dma1_read:slave_read
	wire    [3:0] mm_interconnect_1_video_dma1_read_avalon_dma_control_slave_byteenable;   // mm_interconnect_1:video_dma1_read_avalon_dma_control_slave_byteenable -> video_dma1_read:slave_byteenable
	wire          mm_interconnect_1_video_dma1_read_avalon_dma_control_slave_write;        // mm_interconnect_1:video_dma1_read_avalon_dma_control_slave_write -> video_dma1_read:slave_write
	wire   [31:0] mm_interconnect_1_video_dma1_read_avalon_dma_control_slave_writedata;    // mm_interconnect_1:video_dma1_read_avalon_dma_control_slave_writedata -> video_dma1_read:slave_writedata
	wire   [31:0] mm_interconnect_1_video_dma2_read_avalon_dma_control_slave_readdata;     // video_dma2_read:slave_readdata -> mm_interconnect_1:video_dma2_read_avalon_dma_control_slave_readdata
	wire    [1:0] mm_interconnect_1_video_dma2_read_avalon_dma_control_slave_address;      // mm_interconnect_1:video_dma2_read_avalon_dma_control_slave_address -> video_dma2_read:slave_address
	wire          mm_interconnect_1_video_dma2_read_avalon_dma_control_slave_read;         // mm_interconnect_1:video_dma2_read_avalon_dma_control_slave_read -> video_dma2_read:slave_read
	wire    [3:0] mm_interconnect_1_video_dma2_read_avalon_dma_control_slave_byteenable;   // mm_interconnect_1:video_dma2_read_avalon_dma_control_slave_byteenable -> video_dma2_read:slave_byteenable
	wire          mm_interconnect_1_video_dma2_read_avalon_dma_control_slave_write;        // mm_interconnect_1:video_dma2_read_avalon_dma_control_slave_write -> video_dma2_read:slave_write
	wire   [31:0] mm_interconnect_1_video_dma2_read_avalon_dma_control_slave_writedata;    // mm_interconnect_1:video_dma2_read_avalon_dma_control_slave_writedata -> video_dma2_read:slave_writedata
	wire   [31:0] mm_interconnect_1_alt_vip_vfr_0_avalon_slave_readdata;                   // alt_vip_vfr_0:slave_readdata -> mm_interconnect_1:alt_vip_vfr_0_avalon_slave_readdata
	wire    [4:0] mm_interconnect_1_alt_vip_vfr_0_avalon_slave_address;                    // mm_interconnect_1:alt_vip_vfr_0_avalon_slave_address -> alt_vip_vfr_0:slave_address
	wire          mm_interconnect_1_alt_vip_vfr_0_avalon_slave_read;                       // mm_interconnect_1:alt_vip_vfr_0_avalon_slave_read -> alt_vip_vfr_0:slave_read
	wire          mm_interconnect_1_alt_vip_vfr_0_avalon_slave_write;                      // mm_interconnect_1:alt_vip_vfr_0_avalon_slave_write -> alt_vip_vfr_0:slave_write
	wire   [31:0] mm_interconnect_1_alt_vip_vfr_0_avalon_slave_writedata;                  // mm_interconnect_1:alt_vip_vfr_0_avalon_slave_writedata -> alt_vip_vfr_0:slave_writedata
	wire          pcie_ip_bar2_waitrequest;                                                // mm_interconnect_2:pcie_ip_bar2_waitrequest -> pcie_ip:bar2_waitrequest
	wire   [63:0] pcie_ip_bar2_readdata;                                                   // mm_interconnect_2:pcie_ip_bar2_readdata -> pcie_ip:bar2_readdata
	wire   [31:0] pcie_ip_bar2_address;                                                    // pcie_ip:bar2_address -> mm_interconnect_2:pcie_ip_bar2_address
	wire          pcie_ip_bar2_read;                                                       // pcie_ip:bar2_read -> mm_interconnect_2:pcie_ip_bar2_read
	wire    [7:0] pcie_ip_bar2_byteenable;                                                 // pcie_ip:bar2_byteenable -> mm_interconnect_2:pcie_ip_bar2_byteenable
	wire          pcie_ip_bar2_readdatavalid;                                              // mm_interconnect_2:pcie_ip_bar2_readdatavalid -> pcie_ip:bar2_readdatavalid
	wire          pcie_ip_bar2_write;                                                      // pcie_ip:bar2_write -> mm_interconnect_2:pcie_ip_bar2_write
	wire   [63:0] pcie_ip_bar2_writedata;                                                  // pcie_ip:bar2_writedata -> mm_interconnect_2:pcie_ip_bar2_writedata
	wire    [6:0] pcie_ip_bar2_burstcount;                                                 // pcie_ip:bar2_burstcount -> mm_interconnect_2:pcie_ip_bar2_burstcount
	wire   [31:0] mm_interconnect_2_modular_sgdma_dispatcher_csr_readdata;                 // modular_sgdma_dispatcher:csr_readdata -> mm_interconnect_2:modular_sgdma_dispatcher_CSR_readdata
	wire    [2:0] mm_interconnect_2_modular_sgdma_dispatcher_csr_address;                  // mm_interconnect_2:modular_sgdma_dispatcher_CSR_address -> modular_sgdma_dispatcher:csr_address
	wire          mm_interconnect_2_modular_sgdma_dispatcher_csr_read;                     // mm_interconnect_2:modular_sgdma_dispatcher_CSR_read -> modular_sgdma_dispatcher:csr_read
	wire    [3:0] mm_interconnect_2_modular_sgdma_dispatcher_csr_byteenable;               // mm_interconnect_2:modular_sgdma_dispatcher_CSR_byteenable -> modular_sgdma_dispatcher:csr_byteenable
	wire          mm_interconnect_2_modular_sgdma_dispatcher_csr_write;                    // mm_interconnect_2:modular_sgdma_dispatcher_CSR_write -> modular_sgdma_dispatcher:csr_write
	wire   [31:0] mm_interconnect_2_modular_sgdma_dispatcher_csr_writedata;                // mm_interconnect_2:modular_sgdma_dispatcher_CSR_writedata -> modular_sgdma_dispatcher:csr_writedata
	wire          mm_interconnect_2_modular_sgdma_dispatcher_descriptor_slave_waitrequest; // modular_sgdma_dispatcher:descriptor_waitrequest -> mm_interconnect_2:modular_sgdma_dispatcher_Descriptor_Slave_waitrequest
	wire   [15:0] mm_interconnect_2_modular_sgdma_dispatcher_descriptor_slave_byteenable;  // mm_interconnect_2:modular_sgdma_dispatcher_Descriptor_Slave_byteenable -> modular_sgdma_dispatcher:descriptor_byteenable
	wire          mm_interconnect_2_modular_sgdma_dispatcher_descriptor_slave_write;       // mm_interconnect_2:modular_sgdma_dispatcher_Descriptor_Slave_write -> modular_sgdma_dispatcher:descriptor_write
	wire  [127:0] mm_interconnect_2_modular_sgdma_dispatcher_descriptor_slave_writedata;   // mm_interconnect_2:modular_sgdma_dispatcher_Descriptor_Slave_writedata -> modular_sgdma_dispatcher:descriptor_writedata
	wire          mm_interconnect_2_pcie_ip_cra_chipselect;                                // mm_interconnect_2:pcie_ip_cra_chipselect -> pcie_ip:cra_chipselect
	wire   [31:0] mm_interconnect_2_pcie_ip_cra_readdata;                                  // pcie_ip:cra_readdata -> mm_interconnect_2:pcie_ip_cra_readdata
	wire          mm_interconnect_2_pcie_ip_cra_waitrequest;                               // pcie_ip:cra_waitrequest -> mm_interconnect_2:pcie_ip_cra_waitrequest
	wire   [11:0] mm_interconnect_2_pcie_ip_cra_address;                                   // mm_interconnect_2:pcie_ip_cra_address -> pcie_ip:cra_address
	wire          mm_interconnect_2_pcie_ip_cra_read;                                      // mm_interconnect_2:pcie_ip_cra_read -> pcie_ip:cra_read
	wire    [3:0] mm_interconnect_2_pcie_ip_cra_byteenable;                                // mm_interconnect_2:pcie_ip_cra_byteenable -> pcie_ip:cra_byteenable
	wire          mm_interconnect_2_pcie_ip_cra_write;                                     // mm_interconnect_2:pcie_ip_cra_write -> pcie_ip:cra_write
	wire   [31:0] mm_interconnect_2_pcie_ip_cra_writedata;                                 // mm_interconnect_2:pcie_ip_cra_writedata -> pcie_ip:cra_writedata
	wire          irq_mapper_receiver0_irq;                                                // modular_sgdma_dispatcher:csr_irq -> irq_mapper:receiver0_irq
	wire   [15:0] pcie_ip_rxm_irq_irq;                                                     // irq_mapper:sender_irq -> pcie_ip:rxm_irq_irq
	wire          image_fusion_data_source_valid;                                          // image_fusion:source_valid -> avalon_st_adapter:in_0_valid
	wire   [23:0] image_fusion_data_source_data;                                           // image_fusion:source_data -> avalon_st_adapter:in_0_data
	wire          image_fusion_data_source_ready;                                          // avalon_st_adapter:in_0_ready -> image_fusion:source_ready
	wire          image_fusion_data_source_startofpacket;                                  // image_fusion:source_sop -> avalon_st_adapter:in_0_startofpacket
	wire          image_fusion_data_source_endofpacket;                                    // image_fusion:source_eop -> avalon_st_adapter:in_0_endofpacket
	wire          avalon_st_adapter_out_0_valid;                                           // avalon_st_adapter:out_0_valid -> buffer_write:in_valid
	wire   [23:0] avalon_st_adapter_out_0_data;                                            // avalon_st_adapter:out_0_data -> buffer_write:in_data
	wire          avalon_st_adapter_out_0_ready;                                           // buffer_write:in_ready -> avalon_st_adapter:out_0_ready
	wire          avalon_st_adapter_out_0_startofpacket;                                   // avalon_st_adapter:out_0_startofpacket -> buffer_write:in_startofpacket
	wire          avalon_st_adapter_out_0_endofpacket;                                     // avalon_st_adapter:out_0_endofpacket -> buffer_write:in_endofpacket
	wire    [1:0] avalon_st_adapter_out_0_empty;                                           // avalon_st_adapter:out_0_empty -> buffer_write:in_empty
	wire          buffer_write_out_valid;                                                  // buffer_write:out_valid -> avalon_st_adapter_001:in_0_valid
	wire   [23:0] buffer_write_out_data;                                                   // buffer_write:out_data -> avalon_st_adapter_001:in_0_data
	wire          buffer_write_out_ready;                                                  // avalon_st_adapter_001:in_0_ready -> buffer_write:out_ready
	wire          buffer_write_out_startofpacket;                                          // buffer_write:out_startofpacket -> avalon_st_adapter_001:in_0_startofpacket
	wire          buffer_write_out_endofpacket;                                            // buffer_write:out_endofpacket -> avalon_st_adapter_001:in_0_endofpacket
	wire    [1:0] buffer_write_out_empty;                                                  // buffer_write:out_empty -> avalon_st_adapter_001:in_0_empty
	wire          avalon_st_adapter_001_out_0_valid;                                       // avalon_st_adapter_001:out_0_valid -> video_dma_write:stream_valid
	wire   [23:0] avalon_st_adapter_001_out_0_data;                                        // avalon_st_adapter_001:out_0_data -> video_dma_write:stream_data
	wire          avalon_st_adapter_001_out_0_ready;                                       // video_dma_write:stream_ready -> avalon_st_adapter_001:out_0_ready
	wire          avalon_st_adapter_001_out_0_startofpacket;                               // avalon_st_adapter_001:out_0_startofpacket -> video_dma_write:stream_startofpacket
	wire          avalon_st_adapter_001_out_0_endofpacket;                                 // avalon_st_adapter_001:out_0_endofpacket -> video_dma_write:stream_endofpacket
	wire          rst_controller_reset_out_reset;                                          // rst_controller:reset_out -> [alt_vip_itc_0:rst, alt_vip_vfr_0:master_reset, alt_vip_vfr_0:reset, avalon_st_adapter:in_rst_0_reset, avalon_st_adapter_001:in_rst_0_reset, buffer1_read:reset, buffer2_read:reset, buffer_write:reset, image1_padding:reset, image2_padding:reset, image_fusion:reset, mm_interconnect_0:video_dma1_read_reset_reset_bridge_in_reset_reset, mm_interconnect_1:video_dma_write_reset_reset_bridge_in_reset_reset, sdram:reset_n, video_dma1_read:reset, video_dma2_read:reset, video_dma_write:reset]
	wire          pcie_ip_pcie_core_reset_reset;                                           // pcie_ip:pcie_core_reset_reset_n -> [rst_controller:reset_in1, rst_controller_001:reset_in1, rst_controller_002:reset_in0]
	wire          rst_controller_001_reset_out_reset;                                      // rst_controller_001:reset_out -> altpll_qsys:reset
	wire          rst_controller_002_reset_out_reset;                                      // rst_controller_002:reset_out -> [dma_read_master:reset, dma_write_master:reset, irq_mapper:reset, mm_interconnect_0:dma_read_master_Clock_reset_reset_bridge_in_reset_reset, mm_interconnect_1:pcie_ip_bar1_0_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_2:modular_sgdma_dispatcher_clock_reset_reset_bridge_in_reset_reset, modular_sgdma_dispatcher:reset]

	alt_vipitc131_IS2Vid #(
		.NUMBER_OF_COLOUR_PLANES       (3),
		.COLOUR_PLANES_ARE_IN_PARALLEL (1),
		.BPS                           (8),
		.INTERLACED                    (0),
		.H_ACTIVE_PIXELS               (640),
		.V_ACTIVE_LINES                (480),
		.ACCEPT_COLOURS_IN_SEQ         (0),
		.FIFO_DEPTH                    (12800),
		.CLOCKS_ARE_SAME               (0),
		.USE_CONTROL                   (0),
		.NO_OF_MODES                   (1),
		.THRESHOLD                     (12799),
		.STD_WIDTH                     (1),
		.GENERATE_SYNC                 (0),
		.USE_EMBEDDED_SYNCS            (0),
		.AP_LINE                       (0),
		.V_BLANK                       (0),
		.H_BLANK                       (0),
		.H_SYNC_LENGTH                 (96),
		.H_FRONT_PORCH                 (16),
		.H_BACK_PORCH                  (48),
		.V_SYNC_LENGTH                 (2),
		.V_FRONT_PORCH                 (10),
		.V_BACK_PORCH                  (33),
		.F_RISING_EDGE                 (0),
		.F_FALLING_EDGE                (0),
		.FIELD0_V_RISING_EDGE          (0),
		.FIELD0_V_BLANK                (0),
		.FIELD0_V_SYNC_LENGTH          (0),
		.FIELD0_V_FRONT_PORCH          (0),
		.FIELD0_V_BACK_PORCH           (0),
		.ANC_LINE                      (0),
		.FIELD0_ANC_LINE               (0)
	) alt_vip_itc_0 (
		.is_clk        (altpll_qsys_c0_clk),                                  //       is_clk_rst.clk
		.rst           (rst_controller_reset_out_reset),                      // is_clk_rst_reset.reset
		.is_data       (alt_vip_vfr_0_avalon_streaming_source_data),          //              din.data
		.is_valid      (alt_vip_vfr_0_avalon_streaming_source_valid),         //                 .valid
		.is_ready      (alt_vip_vfr_0_avalon_streaming_source_ready),         //                 .ready
		.is_sop        (alt_vip_vfr_0_avalon_streaming_source_startofpacket), //                 .startofpacket
		.is_eop        (alt_vip_vfr_0_avalon_streaming_source_endofpacket),   //                 .endofpacket
		.vid_clk       (alt_vip_itc_0_clocked_video_vid_clk),                 //    clocked_video.export
		.vid_data      (alt_vip_itc_0_clocked_video_vid_data),                //                 .export
		.underflow     (alt_vip_itc_0_clocked_video_underflow),               //                 .export
		.vid_datavalid (alt_vip_itc_0_clocked_video_vid_datavalid),           //                 .export
		.vid_v_sync    (alt_vip_itc_0_clocked_video_vid_v_sync),              //                 .export
		.vid_h_sync    (alt_vip_itc_0_clocked_video_vid_h_sync),              //                 .export
		.vid_f         (alt_vip_itc_0_clocked_video_vid_f),                   //                 .export
		.vid_h         (alt_vip_itc_0_clocked_video_vid_h),                   //                 .export
		.vid_v         (alt_vip_itc_0_clocked_video_vid_v)                    //                 .export
	);

	alt_vipvfr131_vfr #(
		.BITS_PER_PIXEL_PER_COLOR_PLANE (8),
		.NUMBER_OF_CHANNELS_IN_PARALLEL (3),
		.NUMBER_OF_CHANNELS_IN_SEQUENCE (1),
		.MAX_IMAGE_WIDTH                (640),
		.MAX_IMAGE_HEIGHT               (480),
		.MEM_PORT_WIDTH                 (32),
		.RMASTER_FIFO_DEPTH             (1024),
		.RMASTER_BURST_TARGET           (32),
		.CLOCKS_ARE_SEPARATE            (1)
	) alt_vip_vfr_0 (
		.clock                (altpll_qsys_c0_clk),                                     //             clock_reset.clk
		.reset                (rst_controller_reset_out_reset),                         //       clock_reset_reset.reset
		.master_clock         (altpll_qsys_c0_clk),                                     //            clock_master.clk
		.master_reset         (rst_controller_reset_out_reset),                         //      clock_master_reset.reset
		.slave_address        (mm_interconnect_1_alt_vip_vfr_0_avalon_slave_address),   //            avalon_slave.address
		.slave_write          (mm_interconnect_1_alt_vip_vfr_0_avalon_slave_write),     //                        .write
		.slave_writedata      (mm_interconnect_1_alt_vip_vfr_0_avalon_slave_writedata), //                        .writedata
		.slave_read           (mm_interconnect_1_alt_vip_vfr_0_avalon_slave_read),      //                        .read
		.slave_readdata       (mm_interconnect_1_alt_vip_vfr_0_avalon_slave_readdata),  //                        .readdata
		.slave_irq            (),                                                       //        interrupt_sender.irq
		.dout_data            (alt_vip_vfr_0_avalon_streaming_source_data),             // avalon_streaming_source.data
		.dout_valid           (alt_vip_vfr_0_avalon_streaming_source_valid),            //                        .valid
		.dout_ready           (alt_vip_vfr_0_avalon_streaming_source_ready),            //                        .ready
		.dout_startofpacket   (alt_vip_vfr_0_avalon_streaming_source_startofpacket),    //                        .startofpacket
		.dout_endofpacket     (alt_vip_vfr_0_avalon_streaming_source_endofpacket),      //                        .endofpacket
		.master_address       (alt_vip_vfr_0_avalon_master_address),                    //           avalon_master.address
		.master_burstcount    (alt_vip_vfr_0_avalon_master_burstcount),                 //                        .burstcount
		.master_readdata      (alt_vip_vfr_0_avalon_master_readdata),                   //                        .readdata
		.master_read          (alt_vip_vfr_0_avalon_master_read),                       //                        .read
		.master_readdatavalid (alt_vip_vfr_0_avalon_master_readdatavalid),              //                        .readdatavalid
		.master_waitrequest   (alt_vip_vfr_0_avalon_master_waitrequest)                 //                        .waitrequest
	);

	de2i_150_qsys_altpll_qsys altpll_qsys (
		.clk                (clk_clk),                            //       inclk_interface.clk
		.reset              (rst_controller_001_reset_out_reset), // inclk_interface_reset.reset
		.read               (),                                   //             pll_slave.read
		.write              (),                                   //                      .write
		.address            (),                                   //                      .address
		.readdata           (),                                   //                      .readdata
		.writedata          (),                                   //                      .writedata
		.c0                 (altpll_qsys_c0_clk),                 //                    c0.clk
		.c1                 (altpll_sdram_clk),                   //                    c1.clk
		.c2                 (altpll_vga_clk),                     //                    c2.clk
		.c3                 (altpll_qsys_c3_clk),                 //                    c3.clk
		.c4                 (),                                   //                    c4.clk
		.areset             (),                                   //        areset_conduit.export
		.locked             (),                                   //        locked_conduit.export
		.scandone           (),                                   //           (terminated)
		.scandataout        (),                                   //           (terminated)
		.phasedone          (),                                   //           (terminated)
		.phasecounterselect (4'b0000),                            //           (terminated)
		.phaseupdown        (1'b0),                               //           (terminated)
		.phasestep          (1'b0),                               //           (terminated)
		.scanclk            (1'b0),                               //           (terminated)
		.scanclkena         (1'b0),                               //           (terminated)
		.scandata           (1'b0),                               //           (terminated)
		.configupdate       (1'b0)                                //           (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (8),
		.FIFO_DEPTH          (16384),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (3),
		.USE_MEMORY_BLOCKS   (1),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) buffer1_read (
		.clk               (altpll_qsys_c0_clk),                                //       clk.clk
		.reset             (rst_controller_reset_out_reset),                    // clk_reset.reset
		.in_data           (video_dma1_read_avalon_pixel_source_data),          //        in.data
		.in_valid          (video_dma1_read_avalon_pixel_source_valid),         //          .valid
		.in_ready          (video_dma1_read_avalon_pixel_source_ready),         //          .ready
		.in_startofpacket  (video_dma1_read_avalon_pixel_source_startofpacket), //          .startofpacket
		.in_endofpacket    (video_dma1_read_avalon_pixel_source_endofpacket),   //          .endofpacket
		.out_data          (buffer1_read_out_data),                             //       out.data
		.out_valid         (buffer1_read_out_valid),                            //          .valid
		.out_ready         (buffer1_read_out_ready),                            //          .ready
		.out_startofpacket (buffer1_read_out_startofpacket),                    //          .startofpacket
		.out_endofpacket   (buffer1_read_out_endofpacket),                      //          .endofpacket
		.csr_address       (2'b00),                                             // (terminated)
		.csr_read          (1'b0),                                              // (terminated)
		.csr_write         (1'b0),                                              // (terminated)
		.csr_readdata      (),                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),              // (terminated)
		.almost_full_data  (),                                                  // (terminated)
		.almost_empty_data (),                                                  // (terminated)
		.in_empty          (1'b0),                                              // (terminated)
		.out_empty         (),                                                  // (terminated)
		.in_error          (1'b0),                                              // (terminated)
		.out_error         (),                                                  // (terminated)
		.in_channel        (1'b0),                                              // (terminated)
		.out_channel       ()                                                   // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (8),
		.FIFO_DEPTH          (16384),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (3),
		.USE_MEMORY_BLOCKS   (1),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) buffer2_read (
		.clk               (altpll_qsys_c0_clk),                                //       clk.clk
		.reset             (rst_controller_reset_out_reset),                    // clk_reset.reset
		.in_data           (video_dma2_read_avalon_pixel_source_data),          //        in.data
		.in_valid          (video_dma2_read_avalon_pixel_source_valid),         //          .valid
		.in_ready          (video_dma2_read_avalon_pixel_source_ready),         //          .ready
		.in_startofpacket  (video_dma2_read_avalon_pixel_source_startofpacket), //          .startofpacket
		.in_endofpacket    (video_dma2_read_avalon_pixel_source_endofpacket),   //          .endofpacket
		.out_data          (buffer2_read_out_data),                             //       out.data
		.out_valid         (buffer2_read_out_valid),                            //          .valid
		.out_ready         (buffer2_read_out_ready),                            //          .ready
		.out_startofpacket (buffer2_read_out_startofpacket),                    //          .startofpacket
		.out_endofpacket   (buffer2_read_out_endofpacket),                      //          .endofpacket
		.csr_address       (2'b00),                                             // (terminated)
		.csr_read          (1'b0),                                              // (terminated)
		.csr_write         (1'b0),                                              // (terminated)
		.csr_readdata      (),                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),              // (terminated)
		.almost_full_data  (),                                                  // (terminated)
		.almost_empty_data (),                                                  // (terminated)
		.in_empty          (1'b0),                                              // (terminated)
		.out_empty         (),                                                  // (terminated)
		.in_error          (1'b0),                                              // (terminated)
		.out_error         (),                                                  // (terminated)
		.in_channel        (1'b0),                                              // (terminated)
		.out_channel       ()                                                   // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (3),
		.BITS_PER_SYMBOL     (8),
		.FIFO_DEPTH          (16384),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (3),
		.USE_MEMORY_BLOCKS   (1),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) buffer_write (
		.clk               (altpll_qsys_c0_clk),                    //       clk.clk
		.reset             (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_data           (avalon_st_adapter_out_0_data),          //        in.data
		.in_valid          (avalon_st_adapter_out_0_valid),         //          .valid
		.in_ready          (avalon_st_adapter_out_0_ready),         //          .ready
		.in_startofpacket  (avalon_st_adapter_out_0_startofpacket), //          .startofpacket
		.in_endofpacket    (avalon_st_adapter_out_0_endofpacket),   //          .endofpacket
		.in_empty          (avalon_st_adapter_out_0_empty),         //          .empty
		.out_data          (buffer_write_out_data),                 //       out.data
		.out_valid         (buffer_write_out_valid),                //          .valid
		.out_ready         (buffer_write_out_ready),                //          .ready
		.out_startofpacket (buffer_write_out_startofpacket),        //          .startofpacket
		.out_endofpacket   (buffer_write_out_endofpacket),          //          .endofpacket
		.out_empty         (buffer_write_out_empty),                //          .empty
		.csr_address       (2'b00),                                 // (terminated)
		.csr_read          (1'b0),                                  // (terminated)
		.csr_write         (1'b0),                                  // (terminated)
		.csr_readdata      (),                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),  // (terminated)
		.almost_full_data  (),                                      // (terminated)
		.almost_empty_data (),                                      // (terminated)
		.in_error          (1'b0),                                  // (terminated)
		.out_error         (),                                      // (terminated)
		.in_channel        (1'b0),                                  // (terminated)
		.out_channel       ()                                       // (terminated)
	);

	read_master #(
		.DATA_WIDTH                (32),
		.LENGTH_WIDTH              (23),
		.FIFO_DEPTH                (4096),
		.STRIDE_ENABLE             (0),
		.BURST_ENABLE              (1),
		.PACKET_ENABLE             (0),
		.ERROR_ENABLE              (0),
		.ERROR_WIDTH               (8),
		.CHANNEL_ENABLE            (0),
		.CHANNEL_WIDTH             (8),
		.BYTE_ENABLE_WIDTH         (4),
		.BYTE_ENABLE_WIDTH_LOG2    (2),
		.ADDRESS_WIDTH             (32),
		.FIFO_DEPTH_LOG2           (12),
		.SYMBOL_WIDTH              (8),
		.NUMBER_OF_SYMBOLS         (4),
		.NUMBER_OF_SYMBOLS_LOG2    (2),
		.MAX_BURST_COUNT_WIDTH     (5),
		.UNALIGNED_ACCESSES_ENABLE (1),
		.ONLY_FULL_ACCESS_ENABLE   (0),
		.BURST_WRAPPING_SUPPORT    (0),
		.PROGRAMMABLE_BURST_ENABLE (0),
		.MAX_BURST_COUNT           (16),
		.FIFO_SPEED_OPTIMIZATION   (1),
		.STRIDE_WIDTH              (1)
	) dma_read_master (
		.clk                  (pcie_ip_pcie_core_clk_clk),                          //            Clock.clk
		.reset                (rst_controller_002_reset_out_reset),                 //      Clock_reset.reset
		.master_address       (dma_read_master_data_read_master_address),           // Data_Read_Master.address
		.master_read          (dma_read_master_data_read_master_read),              //                 .read
		.master_byteenable    (dma_read_master_data_read_master_byteenable),        //                 .byteenable
		.master_readdata      (dma_read_master_data_read_master_readdata),          //                 .readdata
		.master_waitrequest   (dma_read_master_data_read_master_waitrequest),       //                 .waitrequest
		.master_readdatavalid (dma_read_master_data_read_master_readdatavalid),     //                 .readdatavalid
		.master_burstcount    (dma_read_master_data_read_master_burstcount),        //                 .burstcount
		.src_data             (dma_read_master_data_source_data),                   //      Data_Source.data
		.src_valid            (dma_read_master_data_source_valid),                  //                 .valid
		.src_ready            (dma_read_master_data_source_ready),                  //                 .ready
		.snk_command_data     (modular_sgdma_dispatcher_read_command_source_data),  //     Command_Sink.data
		.snk_command_valid    (modular_sgdma_dispatcher_read_command_source_valid), //                 .valid
		.snk_command_ready    (modular_sgdma_dispatcher_read_command_source_ready), //                 .ready
		.src_response_data    (dma_read_master_response_source_data),               //  Response_Source.data
		.src_response_valid   (dma_read_master_response_source_valid),              //                 .valid
		.src_response_ready   (dma_read_master_response_source_ready),              //                 .ready
		.src_sop              (),                                                   //      (terminated)
		.src_eop              (),                                                   //      (terminated)
		.src_empty            (),                                                   //      (terminated)
		.src_error            (),                                                   //      (terminated)
		.src_channel          ()                                                    //      (terminated)
	);

	write_master #(
		.DATA_WIDTH                     (32),
		.LENGTH_WIDTH                   (23),
		.FIFO_DEPTH                     (4096),
		.STRIDE_ENABLE                  (0),
		.BURST_ENABLE                   (1),
		.PACKET_ENABLE                  (0),
		.ERROR_ENABLE                   (0),
		.ERROR_WIDTH                    (8),
		.BYTE_ENABLE_WIDTH              (4),
		.BYTE_ENABLE_WIDTH_LOG2         (2),
		.ADDRESS_WIDTH                  (32),
		.FIFO_DEPTH_LOG2                (12),
		.SYMBOL_WIDTH                   (8),
		.NUMBER_OF_SYMBOLS              (4),
		.NUMBER_OF_SYMBOLS_LOG2         (2),
		.MAX_BURST_COUNT_WIDTH          (5),
		.UNALIGNED_ACCESSES_ENABLE      (1),
		.ONLY_FULL_ACCESS_ENABLE        (0),
		.BURST_WRAPPING_SUPPORT         (0),
		.PROGRAMMABLE_BURST_ENABLE      (0),
		.MAX_BURST_COUNT                (16),
		.FIFO_SPEED_OPTIMIZATION        (1),
		.STRIDE_WIDTH                   (1),
		.ACTUAL_BYTES_TRANSFERRED_WIDTH (32)
	) dma_write_master (
		.clk                (pcie_ip_pcie_core_clk_clk),                           //             Clock.clk
		.reset              (rst_controller_002_reset_out_reset),                  //       Clock_reset.reset
		.master_address     (dma_write_master_data_write_master_address),          // Data_Write_Master.address
		.master_write       (dma_write_master_data_write_master_write),            //                  .write
		.master_byteenable  (dma_write_master_data_write_master_byteenable),       //                  .byteenable
		.master_writedata   (dma_write_master_data_write_master_writedata),        //                  .writedata
		.master_waitrequest (dma_write_master_data_write_master_waitrequest),      //                  .waitrequest
		.master_burstcount  (dma_write_master_data_write_master_burstcount),       //                  .burstcount
		.snk_data           (dma_read_master_data_source_data),                    //         Data_Sink.data
		.snk_valid          (dma_read_master_data_source_valid),                   //                  .valid
		.snk_ready          (dma_read_master_data_source_ready),                   //                  .ready
		.snk_command_data   (modular_sgdma_dispatcher_write_command_source_data),  //      Command_Sink.data
		.snk_command_valid  (modular_sgdma_dispatcher_write_command_source_valid), //                  .valid
		.snk_command_ready  (modular_sgdma_dispatcher_write_command_source_ready), //                  .ready
		.src_response_data  (dma_write_master_response_source_data),               //   Response_Source.data
		.src_response_valid (dma_write_master_response_source_valid),              //                  .valid
		.src_response_ready (dma_write_master_response_source_ready),              //                  .ready
		.snk_sop            (1'b0),                                                //       (terminated)
		.snk_eop            (1'b0),                                                //       (terminated)
		.snk_empty          (2'b00),                                               //       (terminated)
		.snk_error          (8'b00000000)                                          //       (terminated)
	);

	de2i_150_qsys_image1_padding image1_padding (
		.clk                      (altpll_qsys_c0_clk),                                 //                   clk.clk
		.reset                    (rst_controller_reset_out_reset),                     //                 reset.reset
		.stream_in_data           (buffer1_read_out_data),                              //   avalon_clipper_sink.data
		.stream_in_startofpacket  (buffer1_read_out_startofpacket),                     //                      .startofpacket
		.stream_in_endofpacket    (buffer1_read_out_endofpacket),                       //                      .endofpacket
		.stream_in_valid          (buffer1_read_out_valid),                             //                      .valid
		.stream_in_ready          (buffer1_read_out_ready),                             //                      .ready
		.stream_out_ready         (image1_padding_avalon_clipper_source_ready),         // avalon_clipper_source.ready
		.stream_out_data          (image1_padding_avalon_clipper_source_data),          //                      .data
		.stream_out_startofpacket (image1_padding_avalon_clipper_source_startofpacket), //                      .startofpacket
		.stream_out_endofpacket   (image1_padding_avalon_clipper_source_endofpacket),   //                      .endofpacket
		.stream_out_valid         (image1_padding_avalon_clipper_source_valid)          //                      .valid
	);

	de2i_150_qsys_image1_padding image2_padding (
		.clk                      (altpll_qsys_c0_clk),                                 //                   clk.clk
		.reset                    (rst_controller_reset_out_reset),                     //                 reset.reset
		.stream_in_data           (buffer2_read_out_data),                              //   avalon_clipper_sink.data
		.stream_in_startofpacket  (buffer2_read_out_startofpacket),                     //                      .startofpacket
		.stream_in_endofpacket    (buffer2_read_out_endofpacket),                       //                      .endofpacket
		.stream_in_valid          (buffer2_read_out_valid),                             //                      .valid
		.stream_in_ready          (buffer2_read_out_ready),                             //                      .ready
		.stream_out_ready         (image2_padding_avalon_clipper_source_ready),         // avalon_clipper_source.ready
		.stream_out_data          (image2_padding_avalon_clipper_source_data),          //                      .data
		.stream_out_startofpacket (image2_padding_avalon_clipper_source_startofpacket), //                      .startofpacket
		.stream_out_endofpacket   (image2_padding_avalon_clipper_source_endofpacket),   //                      .endofpacket
		.stream_out_valid         (image2_padding_avalon_clipper_source_valid)          //                      .valid
	);

	localedgepreserve image_fusion (
		.reset        (rst_controller_reset_out_reset),                     //       reset.reset
		.Clock        (altpll_qsys_c0_clk),                                 //       clock.clk
		.source_data  (image_fusion_data_source_data),                      // data_source.data
		.source_eop   (image_fusion_data_source_endofpacket),               //            .endofpacket
		.source_ready (image_fusion_data_source_ready),                     //            .ready
		.source_sop   (image_fusion_data_source_startofpacket),             //            .startofpacket
		.source_valid (image_fusion_data_source_valid),                     //            .valid
		.sink2_data   (image2_padding_avalon_clipper_source_data),          //  data2_sink.data
		.sink2_eop    (image2_padding_avalon_clipper_source_endofpacket),   //            .endofpacket
		.sink2_ready  (image2_padding_avalon_clipper_source_ready),         //            .ready
		.sink2_sop    (image2_padding_avalon_clipper_source_startofpacket), //            .startofpacket
		.sink2_valid  (image2_padding_avalon_clipper_source_valid),         //            .valid
		.sink1_data   (image1_padding_avalon_clipper_source_data),          //  data1_sink.data
		.sink1_eop    (image1_padding_avalon_clipper_source_endofpacket),   //            .endofpacket
		.sink1_ready  (image1_padding_avalon_clipper_source_ready),         //            .ready
		.sink1_sop    (image1_padding_avalon_clipper_source_startofpacket), //            .startofpacket
		.sink1_valid  (image1_padding_avalon_clipper_source_valid),         //            .valid
		.switch       (switch_name)                                         //      switch.name
	);

	dispatcher #(
		.MODE                        (0),
		.RESPONSE_PORT               (2),
		.DESCRIPTOR_INTERFACE        (0),
		.DESCRIPTOR_FIFO_DEPTH       (8),
		.ENHANCED_FEATURES           (0),
		.DESCRIPTOR_WIDTH            (128),
		.DESCRIPTOR_BYTEENABLE_WIDTH (16)
	) modular_sgdma_dispatcher (
		.clk                     (pcie_ip_pcie_core_clk_clk),                                                                                                             //                clock.clk
		.reset                   (rst_controller_002_reset_out_reset),                                                                                                    //          clock_reset.reset
		.csr_writedata           (mm_interconnect_2_modular_sgdma_dispatcher_csr_writedata),                                                                              //                  CSR.writedata
		.csr_write               (mm_interconnect_2_modular_sgdma_dispatcher_csr_write),                                                                                  //                     .write
		.csr_byteenable          (mm_interconnect_2_modular_sgdma_dispatcher_csr_byteenable),                                                                             //                     .byteenable
		.csr_readdata            (mm_interconnect_2_modular_sgdma_dispatcher_csr_readdata),                                                                               //                     .readdata
		.csr_read                (mm_interconnect_2_modular_sgdma_dispatcher_csr_read),                                                                                   //                     .read
		.csr_address             (mm_interconnect_2_modular_sgdma_dispatcher_csr_address),                                                                                //                     .address
		.descriptor_write        (mm_interconnect_2_modular_sgdma_dispatcher_descriptor_slave_write),                                                                     //     Descriptor_Slave.write
		.descriptor_waitrequest  (mm_interconnect_2_modular_sgdma_dispatcher_descriptor_slave_waitrequest),                                                               //                     .waitrequest
		.descriptor_writedata    (mm_interconnect_2_modular_sgdma_dispatcher_descriptor_slave_writedata),                                                                 //                     .writedata
		.descriptor_byteenable   (mm_interconnect_2_modular_sgdma_dispatcher_descriptor_slave_byteenable),                                                                //                     .byteenable
		.src_write_master_data   (modular_sgdma_dispatcher_write_command_source_data),                                                                                    // Write_Command_Source.data
		.src_write_master_valid  (modular_sgdma_dispatcher_write_command_source_valid),                                                                                   //                     .valid
		.src_write_master_ready  (modular_sgdma_dispatcher_write_command_source_ready),                                                                                   //                     .ready
		.snk_write_master_data   (dma_write_master_response_source_data),                                                                                                 //  Write_Response_Sink.data
		.snk_write_master_valid  (dma_write_master_response_source_valid),                                                                                                //                     .valid
		.snk_write_master_ready  (dma_write_master_response_source_ready),                                                                                                //                     .ready
		.src_read_master_data    (modular_sgdma_dispatcher_read_command_source_data),                                                                                     //  Read_Command_Source.data
		.src_read_master_valid   (modular_sgdma_dispatcher_read_command_source_valid),                                                                                    //                     .valid
		.src_read_master_ready   (modular_sgdma_dispatcher_read_command_source_ready),                                                                                    //                     .ready
		.snk_read_master_data    (dma_read_master_response_source_data),                                                                                                  //   Read_Response_Sink.data
		.snk_read_master_valid   (dma_read_master_response_source_valid),                                                                                                 //                     .valid
		.snk_read_master_ready   (dma_read_master_response_source_ready),                                                                                                 //                     .ready
		.csr_irq                 (irq_mapper_receiver0_irq),                                                                                                              //              csr_irq.irq
		.src_response_data       (),                                                                                                                                      //          (terminated)
		.src_response_valid      (),                                                                                                                                      //          (terminated)
		.src_response_ready      (1'b0),                                                                                                                                  //          (terminated)
		.snk_descriptor_data     (128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000), //          (terminated)
		.snk_descriptor_valid    (1'b0),                                                                                                                                  //          (terminated)
		.snk_descriptor_ready    (),                                                                                                                                      //          (terminated)
		.mm_response_waitrequest (),                                                                                                                                      //          (terminated)
		.mm_response_byteenable  (4'b0000),                                                                                                                               //          (terminated)
		.mm_response_address     (1'b0),                                                                                                                                  //          (terminated)
		.mm_response_readdata    (),                                                                                                                                      //          (terminated)
		.mm_response_read        (1'b0)                                                                                                                                   //          (terminated)
	);

	de2i_150_qsys_pcie_ip #(
		.p_pcie_hip_type                     ("2"),
		.lane_mask                           (8'b11111110),
		.max_link_width                      (1),
		.millisecond_cycle_count             ("125000"),
		.enable_gen2_core                    ("false"),
		.gen2_lane_rate_mode                 ("false"),
		.no_soft_reset                       ("false"),
		.core_clk_divider                    (2),
		.enable_ch0_pclk_out                 ("true"),
		.core_clk_source                     ("pclk"),
		.CB_P2A_AVALON_ADDR_B0               (0),
		.bar0_size_mask                      (8),
		.bar0_io_space                       ("false"),
		.bar0_64bit_mem_space                ("true"),
		.bar0_prefetchable                   ("true"),
		.CB_P2A_AVALON_ADDR_B1               (0),
		.bar1_size_mask                      (0),
		.bar1_io_space                       ("false"),
		.bar1_64bit_mem_space                ("true"),
		.bar1_prefetchable                   ("false"),
		.CB_P2A_AVALON_ADDR_B2               (0),
		.bar2_size_mask                      (26),
		.bar2_io_space                       ("false"),
		.bar2_64bit_mem_space                ("false"),
		.bar2_prefetchable                   ("false"),
		.CB_P2A_AVALON_ADDR_B3               (0),
		.bar3_size_mask                      (0),
		.bar3_io_space                       ("false"),
		.bar3_64bit_mem_space                ("false"),
		.bar3_prefetchable                   ("false"),
		.CB_P2A_AVALON_ADDR_B4               (0),
		.bar4_size_mask                      (0),
		.bar4_io_space                       ("false"),
		.bar4_64bit_mem_space                ("false"),
		.bar4_prefetchable                   ("false"),
		.CB_P2A_AVALON_ADDR_B5               (0),
		.bar5_size_mask                      (0),
		.bar5_io_space                       ("false"),
		.bar5_64bit_mem_space                ("false"),
		.bar5_prefetchable                   ("false"),
		.vendor_id                           (4466),
		.device_id                           (57345),
		.revision_id                         (1),
		.class_code                          (0),
		.subsystem_vendor_id                 (4466),
		.subsystem_device_id                 (4),
		.port_link_number                    (1),
		.msi_function_count                  (0),
		.enable_msi_64bit_addressing         ("true"),
		.enable_function_msix_support        ("false"),
		.eie_before_nfts_count               (4),
		.enable_completion_timeout_disable   ("false"),
		.completion_timeout                  ("NONE"),
		.enable_adapter_half_rate_mode       ("false"),
		.msix_pba_bir                        (0),
		.msix_pba_offset                     (0),
		.msix_table_bir                      (0),
		.msix_table_offset                   (0),
		.msix_table_size                     (0),
		.use_crc_forwarding                  ("false"),
		.surprise_down_error_support         ("false"),
		.dll_active_report_support           ("false"),
		.bar_io_window_size                  ("32BIT"),
		.bar_prefetchable                    (32),
		.hot_plug_support                    (7'b0000000),
		.no_command_completed                ("true"),
		.slot_power_limit                    (0),
		.slot_power_scale                    (0),
		.slot_number                         (0),
		.enable_slot_register                ("false"),
		.advanced_errors                     ("false"),
		.enable_ecrc_check                   ("false"),
		.enable_ecrc_gen                     ("false"),
		.max_payload_size                    (0),
		.retry_buffer_last_active_address    (255),
		.credit_buffer_allocation_aux        ("ABSOLUTE"),
		.vc0_rx_flow_ctrl_posted_header      (28),
		.vc0_rx_flow_ctrl_posted_data        (198),
		.vc0_rx_flow_ctrl_nonposted_header   (30),
		.vc0_rx_flow_ctrl_nonposted_data     (0),
		.vc0_rx_flow_ctrl_compl_header       (48),
		.vc0_rx_flow_ctrl_compl_data         (256),
		.RX_BUF                              (9),
		.RH_NUM                              (7),
		.G_TAG_NUM0                          (32),
		.endpoint_l0_latency                 (0),
		.endpoint_l1_latency                 (0),
		.enable_l1_aspm                      ("false"),
		.l01_entry_latency                   (31),
		.diffclock_nfts_count                (255),
		.sameclock_nfts_count                (255),
		.l1_exit_latency_sameclock           (7),
		.l1_exit_latency_diffclock           (7),
		.l0_exit_latency_sameclock           (7),
		.l0_exit_latency_diffclock           (7),
		.gen2_diffclock_nfts_count           (255),
		.gen2_sameclock_nfts_count           (255),
		.CG_COMMON_CLOCK_MODE                (1),
		.CB_PCIE_MODE                        (0),
		.AST_LITE                            (0),
		.CB_PCIE_RX_LITE                     (0),
		.CG_RXM_IRQ_NUM                      (16),
		.CG_AVALON_S_ADDR_WIDTH              (20),
		.bypass_tl                           ("false"),
		.CG_IMPL_CRA_AV_SLAVE_PORT           (1),
		.CG_NO_CPL_REORDERING                (0),
		.CG_ENABLE_A2P_INTERRUPT             (0),
		.p_user_msi_enable                   (0),
		.CG_IRQ_BIT_ENA                      (65535),
		.CB_A2P_ADDR_MAP_IS_FIXED            (1),
		.CB_A2P_ADDR_MAP_NUM_ENTRIES         (1),
		.CB_A2P_ADDR_MAP_PASS_THRU_BITS      (31),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_0_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_0_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_1_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_1_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_2_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_2_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_3_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_3_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_4_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_4_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_5_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_5_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_6_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_6_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_7_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_7_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_8_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_8_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_9_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_9_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_10_HIGH (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_10_LOW  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_11_HIGH (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_11_LOW  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_12_HIGH (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_12_LOW  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_13_HIGH (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_13_LOW  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_14_HIGH (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_14_LOW  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_15_HIGH (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_15_LOW  (32'b00000000000000000000000000000000),
		.RXM_DATA_WIDTH                      (64),
		.RXM_BEN_WIDTH                       (8),
		.TL_SELECTION                        (1),
		.pcie_mode                           ("SHARED_MODE"),
		.single_rx_detect                    (1),
		.enable_coreclk_out_half_rate        ("false"),
		.low_priority_vc                     (0),
		.link_width                          (1),
		.cyclone4                            (1)
	) pcie_ip (
		.pcie_core_clk_clk                  (pcie_ip_pcie_core_clk_clk),                   //      pcie_core_clk.clk
		.pcie_core_reset_reset_n            (pcie_ip_pcie_core_reset_reset),               //    pcie_core_reset.reset_n
		.cal_blk_clk_clk                    (altpll_qsys_c3_clk),                          //        cal_blk_clk.clk
		.txs_address                        (mm_interconnect_0_pcie_ip_txs_address),       //                txs.address
		.txs_chipselect                     (mm_interconnect_0_pcie_ip_txs_chipselect),    //                   .chipselect
		.txs_byteenable                     (mm_interconnect_0_pcie_ip_txs_byteenable),    //                   .byteenable
		.txs_readdata                       (mm_interconnect_0_pcie_ip_txs_readdata),      //                   .readdata
		.txs_writedata                      (mm_interconnect_0_pcie_ip_txs_writedata),     //                   .writedata
		.txs_read                           (mm_interconnect_0_pcie_ip_txs_read),          //                   .read
		.txs_write                          (mm_interconnect_0_pcie_ip_txs_write),         //                   .write
		.txs_burstcount                     (mm_interconnect_0_pcie_ip_txs_burstcount),    //                   .burstcount
		.txs_readdatavalid                  (mm_interconnect_0_pcie_ip_txs_readdatavalid), //                   .readdatavalid
		.txs_waitrequest                    (mm_interconnect_0_pcie_ip_txs_waitrequest),   //                   .waitrequest
		.refclk_export                      (pcie_ip_refclk_export),                       //             refclk.export
		.test_in_test_in                    (pcie_ip_test_in_test_in),                     //            test_in.test_in
		.pcie_rstn_export                   (pcie_ip_pcie_rstn_export),                    //          pcie_rstn.export
		.clocks_sim_clk250_export           (pcie_ip_clocks_sim_clk250_export),            //         clocks_sim.clk250_export
		.clocks_sim_clk500_export           (pcie_ip_clocks_sim_clk500_export),            //                   .clk500_export
		.clocks_sim_clk125_export           (pcie_ip_clocks_sim_clk125_export),            //                   .clk125_export
		.reconfig_busy_busy_altgxb_reconfig (pcie_ip_reconfig_busy_busy_altgxb_reconfig),  //      reconfig_busy.busy_altgxb_reconfig
		.pipe_ext_pipe_mode                 (pcie_ip_pipe_ext_pipe_mode),                  //           pipe_ext.pipe_mode
		.pipe_ext_phystatus_ext             (pcie_ip_pipe_ext_phystatus_ext),              //                   .phystatus_ext
		.pipe_ext_rate_ext                  (pcie_ip_pipe_ext_rate_ext),                   //                   .rate_ext
		.pipe_ext_powerdown_ext             (pcie_ip_pipe_ext_powerdown_ext),              //                   .powerdown_ext
		.pipe_ext_txdetectrx_ext            (pcie_ip_pipe_ext_txdetectrx_ext),             //                   .txdetectrx_ext
		.pipe_ext_rxelecidle0_ext           (pcie_ip_pipe_ext_rxelecidle0_ext),            //                   .rxelecidle0_ext
		.pipe_ext_rxdata0_ext               (pcie_ip_pipe_ext_rxdata0_ext),                //                   .rxdata0_ext
		.pipe_ext_rxstatus0_ext             (pcie_ip_pipe_ext_rxstatus0_ext),              //                   .rxstatus0_ext
		.pipe_ext_rxvalid0_ext              (pcie_ip_pipe_ext_rxvalid0_ext),               //                   .rxvalid0_ext
		.pipe_ext_rxdatak0_ext              (pcie_ip_pipe_ext_rxdatak0_ext),               //                   .rxdatak0_ext
		.pipe_ext_txdata0_ext               (pcie_ip_pipe_ext_txdata0_ext),                //                   .txdata0_ext
		.pipe_ext_txdatak0_ext              (pcie_ip_pipe_ext_txdatak0_ext),               //                   .txdatak0_ext
		.pipe_ext_rxpolarity0_ext           (pcie_ip_pipe_ext_rxpolarity0_ext),            //                   .rxpolarity0_ext
		.pipe_ext_txcompl0_ext              (pcie_ip_pipe_ext_txcompl0_ext),               //                   .txcompl0_ext
		.pipe_ext_txelecidle0_ext           (pcie_ip_pipe_ext_txelecidle0_ext),            //                   .txelecidle0_ext
		.powerdown_pll_powerdown            (),                                            //          powerdown.pll_powerdown
		.powerdown_gxb_powerdown            (),                                            //                   .gxb_powerdown
		.bar1_0_address                     (pcie_ip_bar1_0_address),                      //             bar1_0.address
		.bar1_0_read                        (pcie_ip_bar1_0_read),                         //                   .read
		.bar1_0_waitrequest                 (pcie_ip_bar1_0_waitrequest),                  //                   .waitrequest
		.bar1_0_write                       (pcie_ip_bar1_0_write),                        //                   .write
		.bar1_0_readdatavalid               (pcie_ip_bar1_0_readdatavalid),                //                   .readdatavalid
		.bar1_0_readdata                    (pcie_ip_bar1_0_readdata),                     //                   .readdata
		.bar1_0_writedata                   (pcie_ip_bar1_0_writedata),                    //                   .writedata
		.bar1_0_burstcount                  (pcie_ip_bar1_0_burstcount),                   //                   .burstcount
		.bar1_0_byteenable                  (pcie_ip_bar1_0_byteenable),                   //                   .byteenable
		.bar2_address                       (pcie_ip_bar2_address),                        //               bar2.address
		.bar2_read                          (pcie_ip_bar2_read),                           //                   .read
		.bar2_waitrequest                   (pcie_ip_bar2_waitrequest),                    //                   .waitrequest
		.bar2_write                         (pcie_ip_bar2_write),                          //                   .write
		.bar2_readdatavalid                 (pcie_ip_bar2_readdatavalid),                  //                   .readdatavalid
		.bar2_readdata                      (pcie_ip_bar2_readdata),                       //                   .readdata
		.bar2_writedata                     (pcie_ip_bar2_writedata),                      //                   .writedata
		.bar2_burstcount                    (pcie_ip_bar2_burstcount),                     //                   .burstcount
		.bar2_byteenable                    (pcie_ip_bar2_byteenable),                     //                   .byteenable
		.cra_chipselect                     (mm_interconnect_2_pcie_ip_cra_chipselect),    //                cra.chipselect
		.cra_address                        (mm_interconnect_2_pcie_ip_cra_address),       //                   .address
		.cra_byteenable                     (mm_interconnect_2_pcie_ip_cra_byteenable),    //                   .byteenable
		.cra_read                           (mm_interconnect_2_pcie_ip_cra_read),          //                   .read
		.cra_readdata                       (mm_interconnect_2_pcie_ip_cra_readdata),      //                   .readdata
		.cra_write                          (mm_interconnect_2_pcie_ip_cra_write),         //                   .write
		.cra_writedata                      (mm_interconnect_2_pcie_ip_cra_writedata),     //                   .writedata
		.cra_waitrequest                    (mm_interconnect_2_pcie_ip_cra_waitrequest),   //                   .waitrequest
		.cra_irq_irq                        (),                                            //            cra_irq.irq
		.rxm_irq_irq                        (pcie_ip_rxm_irq_irq),                         //            rxm_irq.irq
		.rx_in_rx_datain_0                  (pcie_ip_rx_in_rx_datain_0),                   //              rx_in.rx_datain_0
		.tx_out_tx_dataout_0                (pcie_ip_tx_out_tx_dataout_0),                 //             tx_out.tx_dataout_0
		.reconfig_togxb_data                (pcie_ip_reconfig_togxb_data),                 //     reconfig_togxb.data
		.reconfig_gxbclk_clk                (altpll_qsys_c3_clk),                          //    reconfig_gxbclk.clk
		.reconfig_fromgxb_0_data            (pcie_ip_reconfig_fromgxb_0_data),             // reconfig_fromgxb_0.data
		.fixedclk_clk                       (pcie_ip_pcie_core_clk_clk)                    //           fixedclk.clk
	);

	de2i_150_qsys_sdram sdram (
		.clk            (altpll_qsys_c0_clk),                       //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_addr),                               //  wire.export
		.zs_ba          (sdram_ba),                                 //      .export
		.zs_cas_n       (sdram_cas_n),                              //      .export
		.zs_cke         (sdram_cke),                                //      .export
		.zs_cs_n        (sdram_cs_n),                               //      .export
		.zs_dq          (sdram_dq),                                 //      .export
		.zs_dqm         (sdram_dqm),                                //      .export
		.zs_ras_n       (sdram_ras_n),                              //      .export
		.zs_we_n        (sdram_we_n)                                //      .export
	);

	de2i_150_qsys_video_dma1_read video_dma1_read (
		.clk                  (altpll_qsys_c0_clk),                                                    //                      clk.clk
		.reset                (rst_controller_reset_out_reset),                                        //                    reset.reset
		.master_address       (video_dma1_read_avalon_dma_master_address),                             //        avalon_dma_master.address
		.master_waitrequest   (video_dma1_read_avalon_dma_master_waitrequest),                         //                         .waitrequest
		.master_arbiterlock   (video_dma1_read_avalon_dma_master_lock),                                //                         .lock
		.master_read          (video_dma1_read_avalon_dma_master_read),                                //                         .read
		.master_readdata      (video_dma1_read_avalon_dma_master_readdata),                            //                         .readdata
		.master_readdatavalid (video_dma1_read_avalon_dma_master_readdatavalid),                       //                         .readdatavalid
		.slave_address        (mm_interconnect_1_video_dma1_read_avalon_dma_control_slave_address),    // avalon_dma_control_slave.address
		.slave_byteenable     (mm_interconnect_1_video_dma1_read_avalon_dma_control_slave_byteenable), //                         .byteenable
		.slave_read           (mm_interconnect_1_video_dma1_read_avalon_dma_control_slave_read),       //                         .read
		.slave_write          (mm_interconnect_1_video_dma1_read_avalon_dma_control_slave_write),      //                         .write
		.slave_writedata      (mm_interconnect_1_video_dma1_read_avalon_dma_control_slave_writedata),  //                         .writedata
		.slave_readdata       (mm_interconnect_1_video_dma1_read_avalon_dma_control_slave_readdata),   //                         .readdata
		.stream_ready         (video_dma1_read_avalon_pixel_source_ready),                             //      avalon_pixel_source.ready
		.stream_data          (video_dma1_read_avalon_pixel_source_data),                              //                         .data
		.stream_startofpacket (video_dma1_read_avalon_pixel_source_startofpacket),                     //                         .startofpacket
		.stream_endofpacket   (video_dma1_read_avalon_pixel_source_endofpacket),                       //                         .endofpacket
		.stream_valid         (video_dma1_read_avalon_pixel_source_valid)                              //                         .valid
	);

	de2i_150_qsys_video_dma2_read video_dma2_read (
		.clk                  (altpll_qsys_c0_clk),                                                    //                      clk.clk
		.reset                (rst_controller_reset_out_reset),                                        //                    reset.reset
		.master_address       (video_dma2_read_avalon_dma_master_address),                             //        avalon_dma_master.address
		.master_waitrequest   (video_dma2_read_avalon_dma_master_waitrequest),                         //                         .waitrequest
		.master_arbiterlock   (video_dma2_read_avalon_dma_master_lock),                                //                         .lock
		.master_read          (video_dma2_read_avalon_dma_master_read),                                //                         .read
		.master_readdata      (video_dma2_read_avalon_dma_master_readdata),                            //                         .readdata
		.master_readdatavalid (video_dma2_read_avalon_dma_master_readdatavalid),                       //                         .readdatavalid
		.slave_address        (mm_interconnect_1_video_dma2_read_avalon_dma_control_slave_address),    // avalon_dma_control_slave.address
		.slave_byteenable     (mm_interconnect_1_video_dma2_read_avalon_dma_control_slave_byteenable), //                         .byteenable
		.slave_read           (mm_interconnect_1_video_dma2_read_avalon_dma_control_slave_read),       //                         .read
		.slave_write          (mm_interconnect_1_video_dma2_read_avalon_dma_control_slave_write),      //                         .write
		.slave_writedata      (mm_interconnect_1_video_dma2_read_avalon_dma_control_slave_writedata),  //                         .writedata
		.slave_readdata       (mm_interconnect_1_video_dma2_read_avalon_dma_control_slave_readdata),   //                         .readdata
		.stream_ready         (video_dma2_read_avalon_pixel_source_ready),                             //      avalon_pixel_source.ready
		.stream_data          (video_dma2_read_avalon_pixel_source_data),                              //                         .data
		.stream_startofpacket (video_dma2_read_avalon_pixel_source_startofpacket),                     //                         .startofpacket
		.stream_endofpacket   (video_dma2_read_avalon_pixel_source_endofpacket),                       //                         .endofpacket
		.stream_valid         (video_dma2_read_avalon_pixel_source_valid)                              //                         .valid
	);

	de2i_150_qsys_video_dma_write video_dma_write (
		.clk                  (altpll_qsys_c0_clk),                                                    //                      clk.clk
		.reset                (rst_controller_reset_out_reset),                                        //                    reset.reset
		.stream_data          (avalon_st_adapter_001_out_0_data),                                      //          avalon_dma_sink.data
		.stream_startofpacket (avalon_st_adapter_001_out_0_startofpacket),                             //                         .startofpacket
		.stream_endofpacket   (avalon_st_adapter_001_out_0_endofpacket),                               //                         .endofpacket
		.stream_valid         (avalon_st_adapter_001_out_0_valid),                                     //                         .valid
		.stream_ready         (avalon_st_adapter_001_out_0_ready),                                     //                         .ready
		.slave_address        (mm_interconnect_1_video_dma_write_avalon_dma_control_slave_address),    // avalon_dma_control_slave.address
		.slave_byteenable     (mm_interconnect_1_video_dma_write_avalon_dma_control_slave_byteenable), //                         .byteenable
		.slave_read           (mm_interconnect_1_video_dma_write_avalon_dma_control_slave_read),       //                         .read
		.slave_write          (mm_interconnect_1_video_dma_write_avalon_dma_control_slave_write),      //                         .write
		.slave_writedata      (mm_interconnect_1_video_dma_write_avalon_dma_control_slave_writedata),  //                         .writedata
		.slave_readdata       (mm_interconnect_1_video_dma_write_avalon_dma_control_slave_readdata),   //                         .readdata
		.master_address       (video_dma_write_avalon_dma_master_address),                             //        avalon_dma_master.address
		.master_waitrequest   (video_dma_write_avalon_dma_master_waitrequest),                         //                         .waitrequest
		.master_write         (video_dma_write_avalon_dma_master_write),                               //                         .write
		.master_writedata     (video_dma_write_avalon_dma_master_writedata)                            //                         .writedata
	);

	de2i_150_qsys_mm_interconnect_0 mm_interconnect_0 (
		.altpll_qsys_c0_clk                                      (altpll_qsys_c0_clk),                              //                                    altpll_qsys_c0.clk
		.pcie_ip_pcie_core_clk_clk                               (pcie_ip_pcie_core_clk_clk),                       //                             pcie_ip_pcie_core_clk.clk
		.dma_read_master_Clock_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),              // dma_read_master_Clock_reset_reset_bridge_in_reset.reset
		.video_dma1_read_reset_reset_bridge_in_reset_reset       (rst_controller_reset_out_reset),                  //       video_dma1_read_reset_reset_bridge_in_reset.reset
		.alt_vip_vfr_0_avalon_master_address                     (alt_vip_vfr_0_avalon_master_address),             //                       alt_vip_vfr_0_avalon_master.address
		.alt_vip_vfr_0_avalon_master_waitrequest                 (alt_vip_vfr_0_avalon_master_waitrequest),         //                                                  .waitrequest
		.alt_vip_vfr_0_avalon_master_burstcount                  (alt_vip_vfr_0_avalon_master_burstcount),          //                                                  .burstcount
		.alt_vip_vfr_0_avalon_master_read                        (alt_vip_vfr_0_avalon_master_read),                //                                                  .read
		.alt_vip_vfr_0_avalon_master_readdata                    (alt_vip_vfr_0_avalon_master_readdata),            //                                                  .readdata
		.alt_vip_vfr_0_avalon_master_readdatavalid               (alt_vip_vfr_0_avalon_master_readdatavalid),       //                                                  .readdatavalid
		.dma_read_master_Data_Read_Master_address                (dma_read_master_data_read_master_address),        //                  dma_read_master_Data_Read_Master.address
		.dma_read_master_Data_Read_Master_waitrequest            (dma_read_master_data_read_master_waitrequest),    //                                                  .waitrequest
		.dma_read_master_Data_Read_Master_burstcount             (dma_read_master_data_read_master_burstcount),     //                                                  .burstcount
		.dma_read_master_Data_Read_Master_byteenable             (dma_read_master_data_read_master_byteenable),     //                                                  .byteenable
		.dma_read_master_Data_Read_Master_read                   (dma_read_master_data_read_master_read),           //                                                  .read
		.dma_read_master_Data_Read_Master_readdata               (dma_read_master_data_read_master_readdata),       //                                                  .readdata
		.dma_read_master_Data_Read_Master_readdatavalid          (dma_read_master_data_read_master_readdatavalid),  //                                                  .readdatavalid
		.dma_write_master_Data_Write_Master_address              (dma_write_master_data_write_master_address),      //                dma_write_master_Data_Write_Master.address
		.dma_write_master_Data_Write_Master_waitrequest          (dma_write_master_data_write_master_waitrequest),  //                                                  .waitrequest
		.dma_write_master_Data_Write_Master_burstcount           (dma_write_master_data_write_master_burstcount),   //                                                  .burstcount
		.dma_write_master_Data_Write_Master_byteenable           (dma_write_master_data_write_master_byteenable),   //                                                  .byteenable
		.dma_write_master_Data_Write_Master_write                (dma_write_master_data_write_master_write),        //                                                  .write
		.dma_write_master_Data_Write_Master_writedata            (dma_write_master_data_write_master_writedata),    //                                                  .writedata
		.video_dma1_read_avalon_dma_master_address               (video_dma1_read_avalon_dma_master_address),       //                 video_dma1_read_avalon_dma_master.address
		.video_dma1_read_avalon_dma_master_waitrequest           (video_dma1_read_avalon_dma_master_waitrequest),   //                                                  .waitrequest
		.video_dma1_read_avalon_dma_master_read                  (video_dma1_read_avalon_dma_master_read),          //                                                  .read
		.video_dma1_read_avalon_dma_master_readdata              (video_dma1_read_avalon_dma_master_readdata),      //                                                  .readdata
		.video_dma1_read_avalon_dma_master_readdatavalid         (video_dma1_read_avalon_dma_master_readdatavalid), //                                                  .readdatavalid
		.video_dma1_read_avalon_dma_master_lock                  (video_dma1_read_avalon_dma_master_lock),          //                                                  .lock
		.video_dma2_read_avalon_dma_master_address               (video_dma2_read_avalon_dma_master_address),       //                 video_dma2_read_avalon_dma_master.address
		.video_dma2_read_avalon_dma_master_waitrequest           (video_dma2_read_avalon_dma_master_waitrequest),   //                                                  .waitrequest
		.video_dma2_read_avalon_dma_master_read                  (video_dma2_read_avalon_dma_master_read),          //                                                  .read
		.video_dma2_read_avalon_dma_master_readdata              (video_dma2_read_avalon_dma_master_readdata),      //                                                  .readdata
		.video_dma2_read_avalon_dma_master_readdatavalid         (video_dma2_read_avalon_dma_master_readdatavalid), //                                                  .readdatavalid
		.video_dma2_read_avalon_dma_master_lock                  (video_dma2_read_avalon_dma_master_lock),          //                                                  .lock
		.video_dma_write_avalon_dma_master_address               (video_dma_write_avalon_dma_master_address),       //                 video_dma_write_avalon_dma_master.address
		.video_dma_write_avalon_dma_master_waitrequest           (video_dma_write_avalon_dma_master_waitrequest),   //                                                  .waitrequest
		.video_dma_write_avalon_dma_master_write                 (video_dma_write_avalon_dma_master_write),         //                                                  .write
		.video_dma_write_avalon_dma_master_writedata             (video_dma_write_avalon_dma_master_writedata),     //                                                  .writedata
		.pcie_ip_txs_address                                     (mm_interconnect_0_pcie_ip_txs_address),           //                                       pcie_ip_txs.address
		.pcie_ip_txs_write                                       (mm_interconnect_0_pcie_ip_txs_write),             //                                                  .write
		.pcie_ip_txs_read                                        (mm_interconnect_0_pcie_ip_txs_read),              //                                                  .read
		.pcie_ip_txs_readdata                                    (mm_interconnect_0_pcie_ip_txs_readdata),          //                                                  .readdata
		.pcie_ip_txs_writedata                                   (mm_interconnect_0_pcie_ip_txs_writedata),         //                                                  .writedata
		.pcie_ip_txs_burstcount                                  (mm_interconnect_0_pcie_ip_txs_burstcount),        //                                                  .burstcount
		.pcie_ip_txs_byteenable                                  (mm_interconnect_0_pcie_ip_txs_byteenable),        //                                                  .byteenable
		.pcie_ip_txs_readdatavalid                               (mm_interconnect_0_pcie_ip_txs_readdatavalid),     //                                                  .readdatavalid
		.pcie_ip_txs_waitrequest                                 (mm_interconnect_0_pcie_ip_txs_waitrequest),       //                                                  .waitrequest
		.pcie_ip_txs_chipselect                                  (mm_interconnect_0_pcie_ip_txs_chipselect),        //                                                  .chipselect
		.sdram_s1_address                                        (mm_interconnect_0_sdram_s1_address),              //                                          sdram_s1.address
		.sdram_s1_write                                          (mm_interconnect_0_sdram_s1_write),                //                                                  .write
		.sdram_s1_read                                           (mm_interconnect_0_sdram_s1_read),                 //                                                  .read
		.sdram_s1_readdata                                       (mm_interconnect_0_sdram_s1_readdata),             //                                                  .readdata
		.sdram_s1_writedata                                      (mm_interconnect_0_sdram_s1_writedata),            //                                                  .writedata
		.sdram_s1_byteenable                                     (mm_interconnect_0_sdram_s1_byteenable),           //                                                  .byteenable
		.sdram_s1_readdatavalid                                  (mm_interconnect_0_sdram_s1_readdatavalid),        //                                                  .readdatavalid
		.sdram_s1_waitrequest                                    (mm_interconnect_0_sdram_s1_waitrequest),          //                                                  .waitrequest
		.sdram_s1_chipselect                                     (mm_interconnect_0_sdram_s1_chipselect)            //                                                  .chipselect
	);

	de2i_150_qsys_mm_interconnect_1 mm_interconnect_1 (
		.altpll_qsys_c0_clk                                          (altpll_qsys_c0_clk),                                                    //                                        altpll_qsys_c0.clk
		.pcie_ip_pcie_core_clk_clk                                   (pcie_ip_pcie_core_clk_clk),                                             //                                 pcie_ip_pcie_core_clk.clk
		.pcie_ip_bar1_0_translator_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                                    // pcie_ip_bar1_0_translator_reset_reset_bridge_in_reset.reset
		.video_dma_write_reset_reset_bridge_in_reset_reset           (rst_controller_reset_out_reset),                                        //           video_dma_write_reset_reset_bridge_in_reset.reset
		.pcie_ip_bar1_0_address                                      (pcie_ip_bar1_0_address),                                                //                                        pcie_ip_bar1_0.address
		.pcie_ip_bar1_0_waitrequest                                  (pcie_ip_bar1_0_waitrequest),                                            //                                                      .waitrequest
		.pcie_ip_bar1_0_burstcount                                   (pcie_ip_bar1_0_burstcount),                                             //                                                      .burstcount
		.pcie_ip_bar1_0_byteenable                                   (pcie_ip_bar1_0_byteenable),                                             //                                                      .byteenable
		.pcie_ip_bar1_0_read                                         (pcie_ip_bar1_0_read),                                                   //                                                      .read
		.pcie_ip_bar1_0_readdata                                     (pcie_ip_bar1_0_readdata),                                               //                                                      .readdata
		.pcie_ip_bar1_0_readdatavalid                                (pcie_ip_bar1_0_readdatavalid),                                          //                                                      .readdatavalid
		.pcie_ip_bar1_0_write                                        (pcie_ip_bar1_0_write),                                                  //                                                      .write
		.pcie_ip_bar1_0_writedata                                    (pcie_ip_bar1_0_writedata),                                              //                                                      .writedata
		.alt_vip_vfr_0_avalon_slave_address                          (mm_interconnect_1_alt_vip_vfr_0_avalon_slave_address),                  //                            alt_vip_vfr_0_avalon_slave.address
		.alt_vip_vfr_0_avalon_slave_write                            (mm_interconnect_1_alt_vip_vfr_0_avalon_slave_write),                    //                                                      .write
		.alt_vip_vfr_0_avalon_slave_read                             (mm_interconnect_1_alt_vip_vfr_0_avalon_slave_read),                     //                                                      .read
		.alt_vip_vfr_0_avalon_slave_readdata                         (mm_interconnect_1_alt_vip_vfr_0_avalon_slave_readdata),                 //                                                      .readdata
		.alt_vip_vfr_0_avalon_slave_writedata                        (mm_interconnect_1_alt_vip_vfr_0_avalon_slave_writedata),                //                                                      .writedata
		.video_dma1_read_avalon_dma_control_slave_address            (mm_interconnect_1_video_dma1_read_avalon_dma_control_slave_address),    //              video_dma1_read_avalon_dma_control_slave.address
		.video_dma1_read_avalon_dma_control_slave_write              (mm_interconnect_1_video_dma1_read_avalon_dma_control_slave_write),      //                                                      .write
		.video_dma1_read_avalon_dma_control_slave_read               (mm_interconnect_1_video_dma1_read_avalon_dma_control_slave_read),       //                                                      .read
		.video_dma1_read_avalon_dma_control_slave_readdata           (mm_interconnect_1_video_dma1_read_avalon_dma_control_slave_readdata),   //                                                      .readdata
		.video_dma1_read_avalon_dma_control_slave_writedata          (mm_interconnect_1_video_dma1_read_avalon_dma_control_slave_writedata),  //                                                      .writedata
		.video_dma1_read_avalon_dma_control_slave_byteenable         (mm_interconnect_1_video_dma1_read_avalon_dma_control_slave_byteenable), //                                                      .byteenable
		.video_dma2_read_avalon_dma_control_slave_address            (mm_interconnect_1_video_dma2_read_avalon_dma_control_slave_address),    //              video_dma2_read_avalon_dma_control_slave.address
		.video_dma2_read_avalon_dma_control_slave_write              (mm_interconnect_1_video_dma2_read_avalon_dma_control_slave_write),      //                                                      .write
		.video_dma2_read_avalon_dma_control_slave_read               (mm_interconnect_1_video_dma2_read_avalon_dma_control_slave_read),       //                                                      .read
		.video_dma2_read_avalon_dma_control_slave_readdata           (mm_interconnect_1_video_dma2_read_avalon_dma_control_slave_readdata),   //                                                      .readdata
		.video_dma2_read_avalon_dma_control_slave_writedata          (mm_interconnect_1_video_dma2_read_avalon_dma_control_slave_writedata),  //                                                      .writedata
		.video_dma2_read_avalon_dma_control_slave_byteenable         (mm_interconnect_1_video_dma2_read_avalon_dma_control_slave_byteenable), //                                                      .byteenable
		.video_dma_write_avalon_dma_control_slave_address            (mm_interconnect_1_video_dma_write_avalon_dma_control_slave_address),    //              video_dma_write_avalon_dma_control_slave.address
		.video_dma_write_avalon_dma_control_slave_write              (mm_interconnect_1_video_dma_write_avalon_dma_control_slave_write),      //                                                      .write
		.video_dma_write_avalon_dma_control_slave_read               (mm_interconnect_1_video_dma_write_avalon_dma_control_slave_read),       //                                                      .read
		.video_dma_write_avalon_dma_control_slave_readdata           (mm_interconnect_1_video_dma_write_avalon_dma_control_slave_readdata),   //                                                      .readdata
		.video_dma_write_avalon_dma_control_slave_writedata          (mm_interconnect_1_video_dma_write_avalon_dma_control_slave_writedata),  //                                                      .writedata
		.video_dma_write_avalon_dma_control_slave_byteenable         (mm_interconnect_1_video_dma_write_avalon_dma_control_slave_byteenable)  //                                                      .byteenable
	);

	de2i_150_qsys_mm_interconnect_2 mm_interconnect_2 (
		.pcie_ip_pcie_core_clk_clk                                        (pcie_ip_pcie_core_clk_clk),                                               //                                      pcie_ip_pcie_core_clk.clk
		.modular_sgdma_dispatcher_clock_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                                      // modular_sgdma_dispatcher_clock_reset_reset_bridge_in_reset.reset
		.pcie_ip_bar2_address                                             (pcie_ip_bar2_address),                                                    //                                               pcie_ip_bar2.address
		.pcie_ip_bar2_waitrequest                                         (pcie_ip_bar2_waitrequest),                                                //                                                           .waitrequest
		.pcie_ip_bar2_burstcount                                          (pcie_ip_bar2_burstcount),                                                 //                                                           .burstcount
		.pcie_ip_bar2_byteenable                                          (pcie_ip_bar2_byteenable),                                                 //                                                           .byteenable
		.pcie_ip_bar2_read                                                (pcie_ip_bar2_read),                                                       //                                                           .read
		.pcie_ip_bar2_readdata                                            (pcie_ip_bar2_readdata),                                                   //                                                           .readdata
		.pcie_ip_bar2_readdatavalid                                       (pcie_ip_bar2_readdatavalid),                                              //                                                           .readdatavalid
		.pcie_ip_bar2_write                                               (pcie_ip_bar2_write),                                                      //                                                           .write
		.pcie_ip_bar2_writedata                                           (pcie_ip_bar2_writedata),                                                  //                                                           .writedata
		.modular_sgdma_dispatcher_CSR_address                             (mm_interconnect_2_modular_sgdma_dispatcher_csr_address),                  //                               modular_sgdma_dispatcher_CSR.address
		.modular_sgdma_dispatcher_CSR_write                               (mm_interconnect_2_modular_sgdma_dispatcher_csr_write),                    //                                                           .write
		.modular_sgdma_dispatcher_CSR_read                                (mm_interconnect_2_modular_sgdma_dispatcher_csr_read),                     //                                                           .read
		.modular_sgdma_dispatcher_CSR_readdata                            (mm_interconnect_2_modular_sgdma_dispatcher_csr_readdata),                 //                                                           .readdata
		.modular_sgdma_dispatcher_CSR_writedata                           (mm_interconnect_2_modular_sgdma_dispatcher_csr_writedata),                //                                                           .writedata
		.modular_sgdma_dispatcher_CSR_byteenable                          (mm_interconnect_2_modular_sgdma_dispatcher_csr_byteenable),               //                                                           .byteenable
		.modular_sgdma_dispatcher_Descriptor_Slave_write                  (mm_interconnect_2_modular_sgdma_dispatcher_descriptor_slave_write),       //                  modular_sgdma_dispatcher_Descriptor_Slave.write
		.modular_sgdma_dispatcher_Descriptor_Slave_writedata              (mm_interconnect_2_modular_sgdma_dispatcher_descriptor_slave_writedata),   //                                                           .writedata
		.modular_sgdma_dispatcher_Descriptor_Slave_byteenable             (mm_interconnect_2_modular_sgdma_dispatcher_descriptor_slave_byteenable),  //                                                           .byteenable
		.modular_sgdma_dispatcher_Descriptor_Slave_waitrequest            (mm_interconnect_2_modular_sgdma_dispatcher_descriptor_slave_waitrequest), //                                                           .waitrequest
		.pcie_ip_cra_address                                              (mm_interconnect_2_pcie_ip_cra_address),                                   //                                                pcie_ip_cra.address
		.pcie_ip_cra_write                                                (mm_interconnect_2_pcie_ip_cra_write),                                     //                                                           .write
		.pcie_ip_cra_read                                                 (mm_interconnect_2_pcie_ip_cra_read),                                      //                                                           .read
		.pcie_ip_cra_readdata                                             (mm_interconnect_2_pcie_ip_cra_readdata),                                  //                                                           .readdata
		.pcie_ip_cra_writedata                                            (mm_interconnect_2_pcie_ip_cra_writedata),                                 //                                                           .writedata
		.pcie_ip_cra_byteenable                                           (mm_interconnect_2_pcie_ip_cra_byteenable),                                //                                                           .byteenable
		.pcie_ip_cra_waitrequest                                          (mm_interconnect_2_pcie_ip_cra_waitrequest),                               //                                                           .waitrequest
		.pcie_ip_cra_chipselect                                           (mm_interconnect_2_pcie_ip_cra_chipselect)                                 //                                                           .chipselect
	);

	de2i_150_qsys_irq_mapper irq_mapper (
		.clk           (pcie_ip_pcie_core_clk_clk),          //       clk.clk
		.reset         (rst_controller_002_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.sender_irq    (pcie_ip_rxm_irq_irq)                 //    sender.irq
	);

	de2i_150_qsys_avalon_st_adapter #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (24),
		.inChannelWidth  (0),
		.inErrorWidth    (0),
		.inUseEmptyPort  (0),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (24),
		.outChannelWidth (0),
		.outErrorWidth   (0),
		.outUseEmptyPort (1),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter (
		.in_clk_0_clk        (altpll_qsys_c0_clk),                     // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_reset_out_reset),         // in_rst_0.reset
		.in_0_data           (image_fusion_data_source_data),          //     in_0.data
		.in_0_valid          (image_fusion_data_source_valid),         //         .valid
		.in_0_ready          (image_fusion_data_source_ready),         //         .ready
		.in_0_startofpacket  (image_fusion_data_source_startofpacket), //         .startofpacket
		.in_0_endofpacket    (image_fusion_data_source_endofpacket),   //         .endofpacket
		.out_0_data          (avalon_st_adapter_out_0_data),           //    out_0.data
		.out_0_valid         (avalon_st_adapter_out_0_valid),          //         .valid
		.out_0_ready         (avalon_st_adapter_out_0_ready),          //         .ready
		.out_0_startofpacket (avalon_st_adapter_out_0_startofpacket),  //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_out_0_endofpacket),    //         .endofpacket
		.out_0_empty         (avalon_st_adapter_out_0_empty)           //         .empty
	);

	de2i_150_qsys_avalon_st_adapter_001 #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (24),
		.inChannelWidth  (0),
		.inErrorWidth    (0),
		.inUseEmptyPort  (1),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (24),
		.outChannelWidth (0),
		.outErrorWidth   (0),
		.outUseEmptyPort (0),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter_001 (
		.in_clk_0_clk        (altpll_qsys_c0_clk),                        // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_reset_out_reset),            // in_rst_0.reset
		.in_0_data           (buffer_write_out_data),                     //     in_0.data
		.in_0_valid          (buffer_write_out_valid),                    //         .valid
		.in_0_ready          (buffer_write_out_ready),                    //         .ready
		.in_0_startofpacket  (buffer_write_out_startofpacket),            //         .startofpacket
		.in_0_endofpacket    (buffer_write_out_endofpacket),              //         .endofpacket
		.in_0_empty          (buffer_write_out_empty),                    //         .empty
		.out_0_data          (avalon_st_adapter_001_out_0_data),          //    out_0.data
		.out_0_valid         (avalon_st_adapter_001_out_0_valid),         //         .valid
		.out_0_ready         (avalon_st_adapter_001_out_0_ready),         //         .ready
		.out_0_startofpacket (avalon_st_adapter_001_out_0_startofpacket), //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_001_out_0_endofpacket)    //         .endofpacket
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.reset_in1      (~pcie_ip_pcie_core_reset_reset), // reset_in1.reset
		.clk            (altpll_qsys_c0_clk),             //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (~pcie_ip_pcie_core_reset_reset),     // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~pcie_ip_pcie_core_reset_reset),     // reset_in0.reset
		.clk            (pcie_ip_pcie_core_clk_clk),          //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
