-- localedgepreserve_GN_localedgepreserve_Fusion_Cal_Weight.vhd

-- Generated using ACDS version 17.1 590

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity localedgepreserve_GN_localedgepreserve_Fusion_Cal_Weight is
	port (
		pixel_in  : in  std_logic_vector(7 downto 0)  := (others => '0'); --  pixel_in.wire
		valid_in  : in  std_logic                     := '0';             --  valid_in.wire
		max_out   : out std_logic_vector(31 downto 0);                    --   max_out.wire
		Clock     : in  std_logic                     := '0';             --     Clock.clk
		reset     : in  std_logic                     := '0';             --          .reset
		addr_in   : in  std_logic_vector(7 downto 0)  := (others => '0'); --   addr_in.wire
		value_out : out std_logic_vector(31 downto 0);                    -- value_out.wire
		eof_in    : in  std_logic                     := '0'              --    eof_in.wire
	);
end entity localedgepreserve_GN_localedgepreserve_Fusion_Cal_Weight;

architecture rtl of localedgepreserve_GN_localedgepreserve_Fusion_Cal_Weight is
	component alt_dspbuilder_clock_GNQFU4PUDH is
		port (
			aclr      : in  std_logic := 'X'; -- reset
			aclr_n    : in  std_logic := 'X'; -- reset_n
			aclr_out  : out std_logic;        -- reset
			clock     : in  std_logic := 'X'; -- clk
			clock_out : out std_logic         -- clk
		);
	end component alt_dspbuilder_clock_GNQFU4PUDH;

	component alt_dspbuilder_port_GN37ALZBS4 is
		port (
			input  : in  std_logic := 'X'; -- wire
			output : out std_logic         -- wire
		);
	end component alt_dspbuilder_port_GN37ALZBS4;

	component alt_dspbuilder_multiplier_GNUSAT2VBO is
		generic (
			aWidth                         : natural := 8;
			Signed                         : natural := 0;
			bWidth                         : natural := 8;
			DEDICATED_MULTIPLIER_CIRCUITRY : string  := "AUTO";
			pipeline                       : integer := 0;
			OutputLsb                      : integer := 0;
			OutputMsb                      : integer := 8
		);
		port (
			aclr      : in  std_logic                                          := 'X';             -- clk
			clock     : in  std_logic                                          := 'X';             -- clk
			dataa     : in  std_logic_vector(aWidth-1 downto 0)                := (others => 'X'); -- wire
			datab     : in  std_logic_vector(bWidth-1 downto 0)                := (others => 'X'); -- wire
			ena       : in  std_logic                                          := 'X';             -- wire
			result    : out std_logic_vector(OutputMsb-OutputLsb+1-1 downto 0);                    -- wire
			user_aclr : in  std_logic                                          := 'X'              -- wire
		);
	end component alt_dspbuilder_multiplier_GNUSAT2VBO;

	component alt_dspbuilder_gnd_GN is
		port (
			output : out std_logic   -- wire
		);
	end component alt_dspbuilder_gnd_GN;

	component alt_dspbuilder_vcc_GN is
		port (
			output : out std_logic   -- wire
		);
	end component alt_dspbuilder_vcc_GN;

	component alt_dspbuilder_cast_GNBBMDRQ7A is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(31 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNBBMDRQ7A;

	component dual_port_ram_sync is
		port (
			clock         : in  std_logic                     := 'X';             -- clk
			data          : in  std_logic_vector(15 downto 0) := (others => 'X'); -- wire
			q             : out std_logic_vector(15 downto 0);                    -- wire
			read_address  : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- wire
			we            : in  std_logic                     := 'X';             -- wire
			write_address : in  std_logic_vector(7 downto 0)  := (others => 'X')  -- wire
		);
	end component dual_port_ram_sync;

	component alt_dspbuilder_multiplexer_GNIM5IEXF4 is
		generic (
			number_inputs          : natural  := 4;
			pipeline               : natural  := 0;
			width                  : positive := 8;
			HDLTYPE                : string   := "STD_LOGIC_VECTOR";
			use_one_hot_select_bus : natural  := 0
		);
		port (
			clock     : in  std_logic                    := 'X';             -- clk
			aclr      : in  std_logic                    := 'X';             -- reset
			sel       : in  std_logic_vector(0 downto 0) := (others => 'X'); -- wire
			result    : out std_logic_vector(8 downto 0);                    -- wire
			ena       : in  std_logic                    := 'X';             -- wire
			user_aclr : in  std_logic                    := 'X';             -- wire
			in0       : in  std_logic_vector(8 downto 0) := (others => 'X'); -- wire
			in1       : in  std_logic_vector(8 downto 0) := (others => 'X')  -- wire
		);
	end component alt_dspbuilder_multiplexer_GNIM5IEXF4;

	component alt_dspbuilder_port_GNA5S4SQDN is
		port (
			input  : in  std_logic_vector(7 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(7 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNA5S4SQDN;

	component dual_port_ram_sync2 is
		port (
			clock         : in  std_logic                     := 'X';             -- clk
			data          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wire
			max           : out std_logic_vector(31 downto 0);                    -- wire
			q             : out std_logic_vector(31 downto 0);                    -- wire
			read_address  : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- wire
			we            : in  std_logic                     := 'X';             -- wire
			write_address : in  std_logic_vector(7 downto 0)  := (others => 'X')  -- wire
		);
	end component dual_port_ram_sync2;

	component alt_dspbuilder_delay_GNTBDM57LR is
		generic (
			ClockPhase : string   := "1";
			BitPattern : string   := "00000001";
			width      : positive := 8;
			use_init   : natural  := 0;
			delay      : positive := 1
		);
		port (
			aclr   : in  std_logic                          := 'X';             -- clk
			clock  : in  std_logic                          := 'X';             -- clk
			ena    : in  std_logic                          := 'X';             -- wire
			input  : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(width-1 downto 0);                    -- wire
			sclr   : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_delay_GNTBDM57LR;

	component alt_dspbuilder_comparator_GN is
		generic (
			Operator  : string  := "Altaeb";
			lpm_width : natural := 8
		);
		port (
			clock  : in  std_logic                              := 'X';             -- clk
			dataa  : in  std_logic_vector(lpm_width-1 downto 0) := (others => 'X'); -- wire
			datab  : in  std_logic_vector(lpm_width-1 downto 0) := (others => 'X'); -- wire
			result : out std_logic;                                                 -- wire
			sclr   : in  std_logic                              := 'X'              -- clk
		);
	end component alt_dspbuilder_comparator_GN;

	component alt_dspbuilder_counter_GNS5ZU7DCJ is
		generic (
			svalue       : string  := "0";
			use_cnt_ena  : string  := "false";
			use_cout     : string  := "false";
			modulus      : integer := 256;
			use_sclr     : string  := "false";
			ndirection   : natural := 1;
			use_usr_aclr : string  := "false";
			width        : natural := 8;
			use_ena      : string  := "false";
			use_sset     : string  := "false";
			use_aload    : string  := "false";
			avalue       : string  := "0";
			use_aset     : string  := "false";
			use_sload    : string  := "false";
			use_cin      : string  := "false"
		);
		port (
			aclr      : in  std_logic                          := 'X';             -- clk
			aload     : in  std_logic                          := 'X';             -- wire
			aset      : in  std_logic                          := 'X';             -- wire
			cin       : in  std_logic                          := 'X';             -- wire
			clock     : in  std_logic                          := 'X';             -- clk
			cnt_ena   : in  std_logic                          := 'X';             -- wire
			cout      : out std_logic;                                             -- wire
			data      : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			direction : in  std_logic                          := 'X';             -- wire
			ena       : in  std_logic                          := 'X';             -- wire
			q         : out std_logic_vector(width-1 downto 0);                    -- wire
			sclr      : in  std_logic                          := 'X';             -- wire
			sload     : in  std_logic                          := 'X';             -- wire
			sset      : in  std_logic                          := 'X';             -- wire
			user_aclr : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_counter_GNS5ZU7DCJ;

	component alt_dspbuilder_pipelined_adder_GNY2JEH574 is
		generic (
			pipeline : integer := 0;
			width    : natural := 0
		);
		port (
			aclr      : in  std_logic                          := 'X';             -- clk
			add_sub   : in  std_logic                          := 'X';             -- wire
			cin       : in  std_logic                          := 'X';             -- wire
			clock     : in  std_logic                          := 'X';             -- clk
			cout      : out std_logic;                                             -- wire
			dataa     : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			datab     : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			ena       : in  std_logic                          := 'X';             -- wire
			result    : out std_logic_vector(width-1 downto 0);                    -- wire
			user_aclr : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_pipelined_adder_GNY2JEH574;

	component alt_dspbuilder_pipelined_adder_GNTWZRTG4I is
		generic (
			pipeline : integer := 0;
			width    : natural := 0
		);
		port (
			aclr      : in  std_logic                          := 'X';             -- clk
			add_sub   : in  std_logic                          := 'X';             -- wire
			cin       : in  std_logic                          := 'X';             -- wire
			clock     : in  std_logic                          := 'X';             -- clk
			cout      : out std_logic;                                             -- wire
			dataa     : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			datab     : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			ena       : in  std_logic                          := 'X';             -- wire
			result    : out std_logic_vector(width-1 downto 0);                    -- wire
			user_aclr : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_pipelined_adder_GNTWZRTG4I;

	component alt_dspbuilder_logical_bit_op_GNA5ZFEL7V is
		generic (
			LogicalOp     : string   := "AltAND";
			number_inputs : positive := 2
		);
		port (
			result : out std_logic;        -- wire
			data0  : in  std_logic := 'X'; -- wire
			data1  : in  std_logic := 'X'  -- wire
		);
	end component alt_dspbuilder_logical_bit_op_GNA5ZFEL7V;

	component alt_dspbuilder_port_GNEPKLLZKY is
		port (
			input  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(31 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNEPKLLZKY;

	component alt_dspbuilder_constant_GNIIAAYRYZ is
		generic (
			BitPattern : string  := "0000";
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(23 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GNIIAAYRYZ;

	component alt_dspbuilder_logical_bit_op_GNKUBZL4TE is
		generic (
			LogicalOp     : string   := "AltAND";
			number_inputs : positive := 2
		);
		port (
			result : out std_logic;        -- wire
			data0  : in  std_logic := 'X'  -- wire
		);
	end component alt_dspbuilder_logical_bit_op_GNKUBZL4TE;

	component alt_dspbuilder_constant_GNTHQFUUUC is
		generic (
			BitPattern : string  := "0000";
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(9 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GNTHQFUUUC;

	component alt_dspbuilder_logical_bit_op_GNUQ2R64DV is
		generic (
			LogicalOp     : string   := "AltAND";
			number_inputs : positive := 2
		);
		port (
			result : out std_logic;        -- wire
			data0  : in  std_logic := 'X'; -- wire
			data1  : in  std_logic := 'X'  -- wire
		);
	end component alt_dspbuilder_logical_bit_op_GNUQ2R64DV;

	component alt_dspbuilder_constant_GNLUER2G5H is
		generic (
			BitPattern : string  := "0000";
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(18 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GNLUER2G5H;

	component alt_dspbuilder_logical_bit_op_GN5A3KLAEC is
		generic (
			LogicalOp     : string   := "AltAND";
			number_inputs : positive := 2
		);
		port (
			result : out std_logic;        -- wire
			data0  : in  std_logic := 'X'; -- wire
			data1  : in  std_logic := 'X'; -- wire
			data2  : in  std_logic := 'X'  -- wire
		);
	end component alt_dspbuilder_logical_bit_op_GN5A3KLAEC;

	component alt_dspbuilder_constant_GNC5NOVIJT is
		generic (
			BitPattern : string  := "0000";
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(7 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GNC5NOVIJT;

	component alt_dspbuilder_constant_GNRSDUIWRP is
		generic (
			BitPattern : string  := "0000";
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(31 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GNRSDUIWRP;

	component alt_dspbuilder_constant_GN5IRMZXKK is
		generic (
			BitPattern : string  := "0000";
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(9 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GN5IRMZXKK;

	component alt_dspbuilder_constant_GNWFCSDEFM is
		generic (
			BitPattern : string  := "0000";
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(15 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GNWFCSDEFM;

	component alt_dspbuilder_multiplexer_GNTG7F5PN7 is
		generic (
			number_inputs          : natural  := 4;
			pipeline               : natural  := 0;
			width                  : positive := 8;
			HDLTYPE                : string   := "STD_LOGIC_VECTOR";
			use_one_hot_select_bus : natural  := 0
		);
		port (
			clock     : in  std_logic                     := 'X';             -- clk
			aclr      : in  std_logic                     := 'X';             -- reset
			sel       : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- wire
			result    : out std_logic_vector(55 downto 0);                    -- wire
			ena       : in  std_logic                     := 'X';             -- wire
			user_aclr : in  std_logic                     := 'X';             -- wire
			in0       : in  std_logic_vector(55 downto 0) := (others => 'X'); -- wire
			in1       : in  std_logic_vector(55 downto 0) := (others => 'X')  -- wire
		);
	end component alt_dspbuilder_multiplexer_GNTG7F5PN7;

	component alt_dspbuilder_multiplexer_GN7X7SG76C is
		generic (
			number_inputs          : natural  := 4;
			pipeline               : natural  := 0;
			width                  : positive := 8;
			HDLTYPE                : string   := "STD_LOGIC_VECTOR";
			use_one_hot_select_bus : natural  := 0
		);
		port (
			clock     : in  std_logic                     := 'X';             -- clk
			aclr      : in  std_logic                     := 'X';             -- reset
			sel       : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- wire
			result    : out std_logic_vector(15 downto 0);                    -- wire
			ena       : in  std_logic                     := 'X';             -- wire
			user_aclr : in  std_logic                     := 'X';             -- wire
			in0       : in  std_logic_vector(15 downto 0) := (others => 'X'); -- wire
			in1       : in  std_logic_vector(15 downto 0) := (others => 'X')  -- wire
		);
	end component alt_dspbuilder_multiplexer_GN7X7SG76C;

	component alt_dspbuilder_multiplexer_GNCMV7Z7A7 is
		generic (
			number_inputs          : natural  := 4;
			pipeline               : natural  := 0;
			width                  : positive := 8;
			HDLTYPE                : string   := "STD_LOGIC_VECTOR";
			use_one_hot_select_bus : natural  := 0
		);
		port (
			clock     : in  std_logic                     := 'X';             -- clk
			aclr      : in  std_logic                     := 'X';             -- reset
			sel       : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- wire
			result    : out std_logic_vector(10 downto 0);                    -- wire
			ena       : in  std_logic                     := 'X';             -- wire
			user_aclr : in  std_logic                     := 'X';             -- wire
			in0       : in  std_logic_vector(10 downto 0) := (others => 'X'); -- wire
			in1       : in  std_logic_vector(10 downto 0) := (others => 'X')  -- wire
		);
	end component alt_dspbuilder_multiplexer_GNCMV7Z7A7;

	component alt_dspbuilder_multiplexer_GNXY3BAFE2 is
		generic (
			number_inputs          : natural  := 4;
			pipeline               : natural  := 0;
			width                  : positive := 8;
			HDLTYPE                : string   := "STD_LOGIC_VECTOR";
			use_one_hot_select_bus : natural  := 0
		);
		port (
			clock     : in  std_logic                     := 'X';             -- clk
			aclr      : in  std_logic                     := 'X';             -- reset
			sel       : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- wire
			result    : out std_logic_vector(10 downto 0);                    -- wire
			ena       : in  std_logic                     := 'X';             -- wire
			user_aclr : in  std_logic                     := 'X';             -- wire
			in0       : in  std_logic_vector(10 downto 0) := (others => 'X'); -- wire
			in1       : in  std_logic_vector(10 downto 0) := (others => 'X')  -- wire
		);
	end component alt_dspbuilder_multiplexer_GNXY3BAFE2;

	component alt_dspbuilder_memdelay_GNSNJI6FHR is
		generic (
			RAMTYPE : string   := "AUTO";
			WIDTH   : positive := 8;
			DELAY   : positive := 1
		);
		port (
			aclr      : in  std_logic                          := 'X';             -- clk
			clock     : in  std_logic                          := 'X';             -- clk
			ena       : in  std_logic                          := 'X';             -- wire
			input     : in  std_logic_vector(WIDTH-1 downto 0) := (others => 'X'); -- wire
			output    : out std_logic_vector(WIDTH-1 downto 0);                    -- wire
			user_aclr : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_memdelay_GNSNJI6FHR;

	component alt_dspbuilder_memdelay_GNMIZKWFE6 is
		generic (
			RAMTYPE : string   := "AUTO";
			WIDTH   : positive := 8;
			DELAY   : positive := 1
		);
		port (
			aclr      : in  std_logic                          := 'X';             -- clk
			clock     : in  std_logic                          := 'X';             -- clk
			ena       : in  std_logic                          := 'X';             -- wire
			input     : in  std_logic_vector(WIDTH-1 downto 0) := (others => 'X'); -- wire
			output    : out std_logic_vector(WIDTH-1 downto 0);                    -- wire
			user_aclr : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_memdelay_GNMIZKWFE6;

	component alt_dspbuilder_memdelay_GN7KC3ZSDB is
		generic (
			RAMTYPE : string   := "AUTO";
			WIDTH   : positive := 8;
			DELAY   : positive := 1
		);
		port (
			aclr      : in  std_logic                          := 'X';             -- clk
			clock     : in  std_logic                          := 'X';             -- clk
			ena       : in  std_logic                          := 'X';             -- wire
			input     : in  std_logic_vector(WIDTH-1 downto 0) := (others => 'X'); -- wire
			output    : out std_logic_vector(WIDTH-1 downto 0);                    -- wire
			user_aclr : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_memdelay_GN7KC3ZSDB;

	component alt_dspbuilder_memdelay_GNXMJOJMJV is
		generic (
			RAMTYPE : string   := "AUTO";
			WIDTH   : positive := 8;
			DELAY   : positive := 1
		);
		port (
			aclr      : in  std_logic                          := 'X';             -- clk
			clock     : in  std_logic                          := 'X';             -- clk
			ena       : in  std_logic                          := 'X';             -- wire
			input     : in  std_logic_vector(WIDTH-1 downto 0) := (others => 'X'); -- wire
			output    : out std_logic_vector(WIDTH-1 downto 0);                    -- wire
			user_aclr : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_memdelay_GNXMJOJMJV;

	component alt_dspbuilder_multiplier_GNXX7E2RLJ is
		generic (
			aWidth                         : natural := 8;
			Signed                         : natural := 0;
			bWidth                         : natural := 8;
			DEDICATED_MULTIPLIER_CIRCUITRY : string  := "AUTO";
			pipeline                       : integer := 0;
			OutputLsb                      : integer := 0;
			OutputMsb                      : integer := 8
		);
		port (
			aclr      : in  std_logic                                          := 'X';             -- clk
			clock     : in  std_logic                                          := 'X';             -- clk
			dataa     : in  std_logic_vector(aWidth-1 downto 0)                := (others => 'X'); -- wire
			datab     : in  std_logic_vector(bWidth-1 downto 0)                := (others => 'X'); -- wire
			ena       : in  std_logic                                          := 'X';             -- wire
			result    : out std_logic_vector(OutputMsb-OutputLsb+1-1 downto 0);                    -- wire
			user_aclr : in  std_logic                                          := 'X'              -- wire
		);
	end component alt_dspbuilder_multiplier_GNXX7E2RLJ;

	component alt_dspbuilder_delay_GNGQ56ZS4N is
		generic (
			ClockPhase : string   := "1";
			BitPattern : string   := "00000001";
			width      : positive := 8;
			use_init   : natural  := 0;
			delay      : positive := 1
		);
		port (
			aclr   : in  std_logic                          := 'X';             -- clk
			clock  : in  std_logic                          := 'X';             -- clk
			ena    : in  std_logic                          := 'X';             -- wire
			input  : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(width-1 downto 0);                    -- wire
			sclr   : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_delay_GNGQ56ZS4N;

	component alt_dspbuilder_delay_GNNQSQIG3K is
		generic (
			ClockPhase : string   := "1";
			BitPattern : string   := "00000001";
			width      : positive := 8;
			use_init   : natural  := 0;
			delay      : positive := 1
		);
		port (
			aclr   : in  std_logic                          := 'X';             -- clk
			clock  : in  std_logic                          := 'X';             -- clk
			ena    : in  std_logic                          := 'X';             -- wire
			input  : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(width-1 downto 0);                    -- wire
			sclr   : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_delay_GNNQSQIG3K;

	component alt_dspbuilder_constant_GNQE5XU76S is
		generic (
			BitPattern : string  := "0000";
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(9 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GNQE5XU76S;

	component alt_dspbuilder_constant_GNCWI5QDAD is
		generic (
			BitPattern : string  := "0000";
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(15 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GNCWI5QDAD;

	component alt_dspbuilder_constant_GNK57PM5EK is
		generic (
			BitPattern : string  := "0000";
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(9 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GNK57PM5EK;

	component alt_dspbuilder_constant_GNSXLT2IGA is
		generic (
			BitPattern : string  := "0000";
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(8 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GNSXLT2IGA;

	component alt_dspbuilder_counter_GNJYRI37NB is
		generic (
			svalue       : string  := "0";
			use_cnt_ena  : string  := "false";
			use_cout     : string  := "false";
			modulus      : integer := 256;
			use_sclr     : string  := "false";
			ndirection   : natural := 1;
			use_usr_aclr : string  := "false";
			width        : natural := 8;
			use_ena      : string  := "false";
			use_sset     : string  := "false";
			use_aload    : string  := "false";
			avalue       : string  := "0";
			use_aset     : string  := "false";
			use_sload    : string  := "false";
			use_cin      : string  := "false"
		);
		port (
			aclr      : in  std_logic                          := 'X';             -- clk
			aload     : in  std_logic                          := 'X';             -- wire
			aset      : in  std_logic                          := 'X';             -- wire
			cin       : in  std_logic                          := 'X';             -- wire
			clock     : in  std_logic                          := 'X';             -- clk
			cnt_ena   : in  std_logic                          := 'X';             -- wire
			cout      : out std_logic;                                             -- wire
			data      : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			direction : in  std_logic                          := 'X';             -- wire
			ena       : in  std_logic                          := 'X';             -- wire
			q         : out std_logic_vector(width-1 downto 0);                    -- wire
			sclr      : in  std_logic                          := 'X';             -- wire
			sload     : in  std_logic                          := 'X';             -- wire
			sset      : in  std_logic                          := 'X';             -- wire
			user_aclr : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_counter_GNJYRI37NB;

	component alt_dspbuilder_multiplexer_GNMRY6PWYH is
		generic (
			number_inputs          : natural  := 4;
			pipeline               : natural  := 0;
			width                  : positive := 8;
			HDLTYPE                : string   := "STD_LOGIC_VECTOR";
			use_one_hot_select_bus : natural  := 0
		);
		port (
			clock     : in  std_logic                     := 'X';             -- clk
			aclr      : in  std_logic                     := 'X';             -- reset
			sel       : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- wire
			result    : out std_logic_vector(16 downto 0);                    -- wire
			ena       : in  std_logic                     := 'X';             -- wire
			user_aclr : in  std_logic                     := 'X';             -- wire
			in0       : in  std_logic_vector(16 downto 0) := (others => 'X'); -- wire
			in1       : in  std_logic_vector(16 downto 0) := (others => 'X')  -- wire
		);
	end component alt_dspbuilder_multiplexer_GNMRY6PWYH;

	component alt_dspbuilder_delay_GNUACQWN66 is
		generic (
			ClockPhase : string   := "1";
			BitPattern : string   := "00000001";
			width      : positive := 8;
			use_init   : natural  := 0;
			delay      : positive := 1
		);
		port (
			aclr   : in  std_logic                          := 'X';             -- clk
			clock  : in  std_logic                          := 'X';             -- clk
			ena    : in  std_logic                          := 'X';             -- wire
			input  : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(width-1 downto 0);                    -- wire
			sclr   : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_delay_GNUACQWN66;

	component alt_dspbuilder_counter_GNPVW56BJJ is
		generic (
			svalue       : string  := "0";
			use_cnt_ena  : string  := "false";
			use_cout     : string  := "false";
			modulus      : integer := 256;
			use_sclr     : string  := "false";
			ndirection   : natural := 1;
			use_usr_aclr : string  := "false";
			width        : natural := 8;
			use_ena      : string  := "false";
			use_sset     : string  := "false";
			use_aload    : string  := "false";
			avalue       : string  := "0";
			use_aset     : string  := "false";
			use_sload    : string  := "false";
			use_cin      : string  := "false"
		);
		port (
			aclr      : in  std_logic                          := 'X';             -- clk
			aload     : in  std_logic                          := 'X';             -- wire
			aset      : in  std_logic                          := 'X';             -- wire
			cin       : in  std_logic                          := 'X';             -- wire
			clock     : in  std_logic                          := 'X';             -- clk
			cnt_ena   : in  std_logic                          := 'X';             -- wire
			cout      : out std_logic;                                             -- wire
			data      : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			direction : in  std_logic                          := 'X';             -- wire
			ena       : in  std_logic                          := 'X';             -- wire
			q         : out std_logic_vector(width-1 downto 0);                    -- wire
			sclr      : in  std_logic                          := 'X';             -- wire
			sload     : in  std_logic                          := 'X';             -- wire
			sset      : in  std_logic                          := 'X';             -- wire
			user_aclr : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_counter_GNPVW56BJJ;

	component alt_dspbuilder_delay_GNQBXYU75H is
		generic (
			ClockPhase : string   := "1";
			BitPattern : string   := "00000001";
			width      : positive := 8;
			use_init   : natural  := 0;
			delay      : positive := 1
		);
		port (
			aclr   : in  std_logic                          := 'X';             -- clk
			clock  : in  std_logic                          := 'X';             -- clk
			ena    : in  std_logic                          := 'X';             -- wire
			input  : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(width-1 downto 0);                    -- wire
			sclr   : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_delay_GNQBXYU75H;

	component alt_dspbuilder_multiplexer_GNWZZP2IFI is
		generic (
			number_inputs          : natural  := 4;
			pipeline               : natural  := 0;
			width                  : positive := 8;
			HDLTYPE                : string   := "STD_LOGIC_VECTOR";
			use_one_hot_select_bus : natural  := 0
		);
		port (
			clock     : in  std_logic                    := 'X';             -- clk
			aclr      : in  std_logic                    := 'X';             -- reset
			sel       : in  std_logic_vector(0 downto 0) := (others => 'X'); -- wire
			result    : out std_logic_vector(9 downto 0);                    -- wire
			ena       : in  std_logic                    := 'X';             -- wire
			user_aclr : in  std_logic                    := 'X';             -- wire
			in0       : in  std_logic_vector(9 downto 0) := (others => 'X'); -- wire
			in1       : in  std_logic_vector(9 downto 0) := (others => 'X')  -- wire
		);
	end component alt_dspbuilder_multiplexer_GNWZZP2IFI;

	component alt_dspbuilder_multiplexer_GNAIWAHV3K is
		generic (
			number_inputs          : natural  := 4;
			pipeline               : natural  := 0;
			width                  : positive := 8;
			HDLTYPE                : string   := "STD_LOGIC_VECTOR";
			use_one_hot_select_bus : natural  := 0
		);
		port (
			clock     : in  std_logic                    := 'X';             -- clk
			aclr      : in  std_logic                    := 'X';             -- reset
			sel       : in  std_logic_vector(0 downto 0) := (others => 'X'); -- wire
			result    : out std_logic_vector(0 downto 0);                    -- wire
			ena       : in  std_logic                    := 'X';             -- wire
			user_aclr : in  std_logic                    := 'X';             -- wire
			in0       : in  std_logic_vector(0 downto 0) := (others => 'X'); -- wire
			in1       : in  std_logic_vector(0 downto 0) := (others => 'X')  -- wire
		);
	end component alt_dspbuilder_multiplexer_GNAIWAHV3K;

	component alt_dspbuilder_cast_GNU3FOKJ6W is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(31 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNU3FOKJ6W;

	component alt_dspbuilder_cast_GNHIWMUP5U is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(31 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNHIWMUP5U;

	component alt_dspbuilder_cast_GNOFO5NIX3 is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(18 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(20 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNOFO5NIX3;

	component alt_dspbuilder_cast_GN6OFM6A6B is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- wire
			output : out std_logic_vector(10 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GN6OFM6A6B;

	component alt_dspbuilder_cast_GN5D52DF5S is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- wire
			output : out std_logic_vector(10 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GN5D52DF5S;

	component alt_dspbuilder_cast_GNAMS3PPNH is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- wire
			output : out std_logic_vector(10 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNAMS3PPNH;

	component alt_dspbuilder_cast_GNSB3OXIQS is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(0 downto 0) := (others => 'X'); -- wire
			output : out std_logic                                        -- wire
		);
	end component alt_dspbuilder_cast_GNSB3OXIQS;

	component alt_dspbuilder_cast_GN5JC4724B is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(19 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(20 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GN5JC4724B;

	component alt_dspbuilder_cast_GNPFJ7B3O7 is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(8 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(9 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNPFJ7B3O7;

	component alt_dspbuilder_cast_GNVKZTMEYW is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(9 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(7 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNVKZTMEYW;

	component alt_dspbuilder_cast_GNBZR5PMEK is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(7 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(7 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNBZR5PMEK;

	component alt_dspbuilder_cast_GNUW2C7J4Q is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(7 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(8 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNUW2C7J4Q;

	component alt_dspbuilder_cast_GNQQ42CR65 is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(15 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNQQ42CR65;

	component alt_dspbuilder_cast_GNSKTJRCBQ is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(8 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(7 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNSKTJRCBQ;

	component alt_dspbuilder_cast_GN46N4UJ5S is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic                    := 'X'; -- wire
			output : out std_logic_vector(0 downto 0)         -- wire
		);
	end component alt_dspbuilder_cast_GN46N4UJ5S;

	component alt_dspbuilder_cast_GNXDXNUGW4 is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(7 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(8 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNXDXNUGW4;

	component alt_dspbuilder_cast_GNRXYRYI2J is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- wire
			output : out std_logic_vector(10 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNRXYRYI2J;

	component alt_dspbuilder_cast_GNBKDIMZSI is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(55 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNBKDIMZSI;

	component alt_dspbuilder_cast_GNNDZ2WJEB is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(7 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(9 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNNDZ2WJEB;

	component alt_dspbuilder_cast_GNOZDXZSET is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(16 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNOZDXZSET;

	component alt_dspbuilder_cast_GNACWQQVMS is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(16 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNACWQQVMS;

	component alt_dspbuilder_cast_GNQ4YFQS5C is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(15 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNQ4YFQS5C;

	component alt_dspbuilder_cast_GNJYJUBV3U is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(10 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(7 downto 0)                      -- wire
		);
	end component alt_dspbuilder_cast_GNJYJUBV3U;

	component alt_dspbuilder_cast_GN5PMHXBFJ is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(16 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(15 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GN5PMHXBFJ;

	component alt_dspbuilder_cast_GNZEACPTPO is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(31 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNZEACPTPO;

	component alt_dspbuilder_cast_GNNQZKMK3E is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(55 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(31 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNNQZKMK3E;

	component alt_dspbuilder_cast_GN5UGBMOKS is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(31 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GN5UGBMOKS;

	component alt_dspbuilder_cast_GNSR6E4BZE is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(55 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNSR6E4BZE;

	component alt_dspbuilder_cast_GNDTOV7QCB is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(10 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(9 downto 0)                      -- wire
		);
	end component alt_dspbuilder_cast_GNDTOV7QCB;

	signal multiplier1user_aclrgnd_output_wire      : std_logic;                     -- Multiplier1user_aclrGND:output -> Multiplier1:user_aclr
	signal multiplier1enavcc_output_wire            : std_logic;                     -- Multiplier1enaVCC:output -> Multiplier1:ena
	signal multiplexeruser_aclrgnd_output_wire      : std_logic;                     -- Multiplexeruser_aclrGND:output -> Multiplexer:user_aclr
	signal multiplexerenavcc_output_wire            : std_logic;                     -- MultiplexerenaVCC:output -> Multiplexer:ena
	signal delaysclrgnd_output_wire                 : std_logic;                     -- DelaysclrGND:output -> Delay:sclr
	signal delayenavcc_output_wire                  : std_logic;                     -- DelayenaVCC:output -> Delay:ena
	signal pipelined_adder2user_aclrgnd_output_wire : std_logic;                     -- Pipelined_Adder2user_aclrGND:output -> Pipelined_Adder2:user_aclr
	signal pipelined_adder2enavcc_output_wire       : std_logic;                     -- Pipelined_Adder2enaVCC:output -> Pipelined_Adder2:ena
	signal pipelined_adder1user_aclrgnd_output_wire : std_logic;                     -- Pipelined_Adder1user_aclrGND:output -> Pipelined_Adder1:user_aclr
	signal pipelined_adder1enavcc_output_wire       : std_logic;                     -- Pipelined_Adder1enaVCC:output -> Pipelined_Adder1:ena
	signal multiplexer3user_aclrgnd_output_wire     : std_logic;                     -- Multiplexer3user_aclrGND:output -> Multiplexer3:user_aclr
	signal multiplexer3enavcc_output_wire           : std_logic;                     -- Multiplexer3enaVCC:output -> Multiplexer3:ena
	signal multiplexer4user_aclrgnd_output_wire     : std_logic;                     -- Multiplexer4user_aclrGND:output -> Multiplexer4:user_aclr
	signal multiplexer4enavcc_output_wire           : std_logic;                     -- Multiplexer4enaVCC:output -> Multiplexer4:ena
	signal multiplexer1user_aclrgnd_output_wire     : std_logic;                     -- Multiplexer1user_aclrGND:output -> Multiplexer1:user_aclr
	signal multiplexer1enavcc_output_wire           : std_logic;                     -- Multiplexer1enaVCC:output -> Multiplexer1:ena
	signal multiplexer2user_aclrgnd_output_wire     : std_logic;                     -- Multiplexer2user_aclrGND:output -> Multiplexer2:user_aclr
	signal multiplexer2enavcc_output_wire           : std_logic;                     -- Multiplexer2enaVCC:output -> Multiplexer2:ena
	signal memory_delay7user_aclrgnd_output_wire    : std_logic;                     -- Memory_Delay7user_aclrGND:output -> Memory_Delay7:user_aclr
	signal memory_delay7enavcc_output_wire          : std_logic;                     -- Memory_Delay7enaVCC:output -> Memory_Delay7:ena
	signal pipelined_adderuser_aclrgnd_output_wire  : std_logic;                     -- Pipelined_Adderuser_aclrGND:output -> Pipelined_Adder:user_aclr
	signal pipelined_adderenavcc_output_wire        : std_logic;                     -- Pipelined_AdderenaVCC:output -> Pipelined_Adder:ena
	signal memory_delay8user_aclrgnd_output_wire    : std_logic;                     -- Memory_Delay8user_aclrGND:output -> Memory_Delay8:user_aclr
	signal memory_delay8enavcc_output_wire          : std_logic;                     -- Memory_Delay8enaVCC:output -> Memory_Delay8:ena
	signal memory_delay5user_aclrgnd_output_wire    : std_logic;                     -- Memory_Delay5user_aclrGND:output -> Memory_Delay5:user_aclr
	signal memory_delay5enavcc_output_wire          : std_logic;                     -- Memory_Delay5enaVCC:output -> Memory_Delay5:ena
	signal memory_delay6user_aclrgnd_output_wire    : std_logic;                     -- Memory_Delay6user_aclrGND:output -> Memory_Delay6:user_aclr
	signal memory_delay6enavcc_output_wire          : std_logic;                     -- Memory_Delay6enaVCC:output -> Memory_Delay6:ena
	signal memory_delay3user_aclrgnd_output_wire    : std_logic;                     -- Memory_Delay3user_aclrGND:output -> Memory_Delay3:user_aclr
	signal memory_delay3enavcc_output_wire          : std_logic;                     -- Memory_Delay3enaVCC:output -> Memory_Delay3:ena
	signal memory_delay4user_aclrgnd_output_wire    : std_logic;                     -- Memory_Delay4user_aclrGND:output -> Memory_Delay4:user_aclr
	signal memory_delay4enavcc_output_wire          : std_logic;                     -- Memory_Delay4enaVCC:output -> Memory_Delay4:ena
	signal memory_delay1user_aclrgnd_output_wire    : std_logic;                     -- Memory_Delay1user_aclrGND:output -> Memory_Delay1:user_aclr
	signal memory_delay1enavcc_output_wire          : std_logic;                     -- Memory_Delay1enaVCC:output -> Memory_Delay1:ena
	signal memory_delay2user_aclrgnd_output_wire    : std_logic;                     -- Memory_Delay2user_aclrGND:output -> Memory_Delay2:user_aclr
	signal memory_delay2enavcc_output_wire          : std_logic;                     -- Memory_Delay2enaVCC:output -> Memory_Delay2:ena
	signal multiplieruser_aclrgnd_output_wire       : std_logic;                     -- Multiplieruser_aclrGND:output -> Multiplier:user_aclr
	signal multiplierenavcc_output_wire             : std_logic;                     -- MultiplierenaVCC:output -> Multiplier:ena
	signal delay2sclrgnd_output_wire                : std_logic;                     -- Delay2sclrGND:output -> Delay2:sclr
	signal delay2enavcc_output_wire                 : std_logic;                     -- Delay2enaVCC:output -> Delay2:ena
	signal delay1sclrgnd_output_wire                : std_logic;                     -- Delay1sclrGND:output -> Delay1:sclr
	signal delay1enavcc_output_wire                 : std_logic;                     -- Delay1enaVCC:output -> Delay1:ena
	signal multiplexer7user_aclrgnd_output_wire     : std_logic;                     -- Multiplexer7user_aclrGND:output -> Multiplexer7:user_aclr
	signal multiplexer7enavcc_output_wire           : std_logic;                     -- Multiplexer7enaVCC:output -> Multiplexer7:ena
	signal delay5sclrgnd_output_wire                : std_logic;                     -- Delay5sclrGND:output -> Delay5:sclr
	signal delay5enavcc_output_wire                 : std_logic;                     -- Delay5enaVCC:output -> Delay5:ena
	signal multiplexer8user_aclrgnd_output_wire     : std_logic;                     -- Multiplexer8user_aclrGND:output -> Multiplexer8:user_aclr
	signal multiplexer8enavcc_output_wire           : std_logic;                     -- Multiplexer8enaVCC:output -> Multiplexer8:ena
	signal delay4sclrgnd_output_wire                : std_logic;                     -- Delay4sclrGND:output -> Delay4:sclr
	signal delay4enavcc_output_wire                 : std_logic;                     -- Delay4enaVCC:output -> Delay4:ena
	signal multiplexer5user_aclrgnd_output_wire     : std_logic;                     -- Multiplexer5user_aclrGND:output -> Multiplexer5:user_aclr
	signal multiplexer5enavcc_output_wire           : std_logic;                     -- Multiplexer5enaVCC:output -> Multiplexer5:ena
	signal multiplexer6user_aclrgnd_output_wire     : std_logic;                     -- Multiplexer6user_aclrGND:output -> Multiplexer6:user_aclr
	signal multiplexer6enavcc_output_wire           : std_logic;                     -- Multiplexer6enaVCC:output -> Multiplexer6:ena
	signal constant5_output_wire                    : std_logic_vector(9 downto 0);  -- Constant5:output -> Comparator1:datab
	signal valid_in_0_output_wire                   : std_logic;                     -- valid_in_0:output -> [Counter:cnt_ena, Logical_Bit_Operator10:data1, Logical_Bit_Operator1:data0, Logical_Bit_Operator8:data1, cast206:input]
	signal delay2_output_wire                       : std_logic_vector(0 downto 0);  -- Delay2:output -> [Delay1:input, Delay4:input, cast190:input, cast200:input]
	signal counter2_q_wire                          : std_logic_vector(9 downto 0);  -- Counter2:q -> [Delay5:input, cast186:input, cast187:input, cast191:input, cast212:input]
	signal logical_bit_operator5_result_wire        : std_logic;                     -- Logical_Bit_Operator5:result -> [Counter2:sclr, Counter3:sclr, Counter:sclr, Logical_Bit_Operator6:data1]
	signal comparator_result_wire                   : std_logic;                     -- Comparator:result -> [Logical_Bit_Operator2:data0, Logical_Bit_Operator7:data0, Logical_Bit_Operator:data0, cast209:input]
	signal logical_bit_operator_result_wire         : std_logic;                     -- Logical_Bit_Operator:result -> Logical_Bit_Operator1:data1
	signal comparator5_result_wire                  : std_logic;                     -- Comparator5:result -> Logical_Bit_Operator10:data0
	signal comparator6_result_wire                  : std_logic;                     -- Comparator6:result -> Logical_Bit_Operator2:data1
	signal logical_bit_operator2_result_wire        : std_logic;                     -- Logical_Bit_Operator2:result -> Counter1:cnt_ena
	signal comparator7_result_wire                  : std_logic;                     -- Comparator7:result -> [Logical_Bit_Operator3:data0, cast216:input, cast217:input, cast219:input]
	signal comparator8_result_wire                  : std_logic;                     -- Comparator8:result -> [Logical_Bit_Operator3:data1, Logical_Bit_Operator4:data0]
	signal logical_bit_operator3_result_wire        : std_logic;                     -- Logical_Bit_Operator3:result -> Counter3:cnt_ena
	signal eof_in_0_output_wire                     : std_logic;                     -- eof_in_0:output -> Logical_Bit_Operator5:data0
	signal logical_bit_operator4_result_wire        : std_logic;                     -- Logical_Bit_Operator4:result -> Logical_Bit_Operator5:data1
	signal logical_bit_operator6_result_wire        : std_logic;                     -- Logical_Bit_Operator6:result -> Counter1:sclr
	signal comparator4_result_wire                  : std_logic;                     -- Comparator4:result -> Logical_Bit_Operator7:data1
	signal comparator2_result_wire                  : std_logic;                     -- Comparator2:result -> Logical_Bit_Operator8:data0
	signal pixel_in_0_output_wire                   : std_logic_vector(7 downto 0);  -- pixel_in_0:output -> [Memory_Delay1:input, Memory_Delay2:input, cast192:input, cast193:input, cast210:input]
	signal memory_delay2_output_wire                : std_logic_vector(7 downto 0);  -- Memory_Delay2:output -> [Memory_Delay4:input, cast202:input]
	signal memory_delay7_output_wire                : std_logic_vector(0 downto 0);  -- Memory_Delay7:output -> [Memory_Delay8:input, cast207:input]
	signal counter1_q_wire                          : std_logic_vector(8 downto 0);  -- Counter1:q -> [Multiplexer:in1, cast184:input, cast194:input]
	signal multiplexer1_result_wire                 : std_logic_vector(10 downto 0); -- Multiplexer1:result -> [Comparator3:dataa, Multiplexer2:in0]
	signal delay1_output_wire                       : std_logic_vector(0 downto 0);  -- Delay1:output -> Multiplexer3:sel
	signal constant13_output_wire                   : std_logic_vector(15 downto 0); -- Constant13:output -> Multiplexer4:in1
	signal multiplexer4_result_wire                 : std_logic_vector(15 downto 0); -- Multiplexer4:result -> [Memory_Delay5:input, cast195:input, cast220:input]
	signal counter3_q_wire                          : std_logic_vector(9 downto 0);  -- Counter3:q -> [Multiplexer5:in1, cast188:input]
	signal delay_output_wire                        : std_logic_vector(0 downto 0);  -- Delay:output -> Multiplexer6:in0
	signal memory_delay3_output_wire                : std_logic_vector(0 downto 0);  -- Memory_Delay3:output -> Multiplexer7:sel
	signal memory_delay6_output_wire                : std_logic_vector(0 downto 0);  -- Memory_Delay6:output -> Multiplexer8:sel
	signal multiplexer8_result_wire                 : std_logic_vector(16 downto 0); -- Multiplexer8:result -> Multiplexer7:in0
	signal constant2_output_wire                    : std_logic_vector(23 downto 0); -- Constant2:output -> Multiplier:datab
	signal multiplier_result_wire                   : std_logic_vector(31 downto 0); -- Multiplier:result -> Binary_Point_Casting:input
	signal constant4_output_wire                    : std_logic_vector(15 downto 0); -- Constant4:output -> Pipelined_Adder:datab
	signal pipelined_adder_result_wire              : std_logic_vector(15 downto 0); -- Pipelined_Adder:result -> Multiplexer4:in0
	signal constant3_output_wire                    : std_logic_vector(9 downto 0);  -- Constant3:output -> Pipelined_Adder2:datab
	signal binary_point_casting1_output_wire        : std_logic_vector(31 downto 0); -- Binary_Point_Casting1:output -> value_out_0:input
	signal binary_point_casting2_output_wire        : std_logic_vector(31 downto 0); -- Binary_Point_Casting2:output -> max_out_0:input
	signal binary_point_casting_output_wire         : std_logic_vector(31 downto 0); -- Binary_Point_Casting:output -> cast174:input
	signal cast174_output_wire                      : std_logic_vector(31 downto 0); -- cast174:output -> Acc_Histogram:data
	signal acc_histogram_q_wire                     : std_logic_vector(31 downto 0); -- Acc_Histogram:q -> cast175:input
	signal cast175_output_wire                      : std_logic_vector(31 downto 0); -- cast175:output -> Binary_Point_Casting1:input
	signal acc_histogram_max_wire                   : std_logic_vector(31 downto 0); -- Acc_Histogram:max -> cast176:input
	signal cast176_output_wire                      : std_logic_vector(31 downto 0); -- cast176:output -> Binary_Point_Casting2:input
	signal constant1_output_wire                    : std_logic_vector(18 downto 0); -- Constant1:output -> cast177:input
	signal cast177_output_wire                      : std_logic_vector(20 downto 0); -- cast177:output -> Comparator:datab
	signal constant11_output_wire                   : std_logic_vector(8 downto 0);  -- Constant11:output -> cast178:input
	signal cast178_output_wire                      : std_logic_vector(10 downto 0); -- cast178:output -> Comparator6:datab
	signal constant12_output_wire                   : std_logic_vector(9 downto 0);  -- Constant12:output -> cast179:input
	signal cast179_output_wire                      : std_logic_vector(10 downto 0); -- cast179:output -> Comparator7:datab
	signal constant14_output_wire                   : std_logic_vector(9 downto 0);  -- Constant14:output -> cast180:input
	signal cast180_output_wire                      : std_logic_vector(10 downto 0); -- cast180:output -> Comparator8:datab
	signal constant7_output_wire                    : std_logic_vector(9 downto 0);  -- Constant7:output -> cast181:input
	signal cast181_output_wire                      : std_logic_vector(10 downto 0); -- cast181:output -> Comparator3:datab
	signal delay4_output_wire                       : std_logic_vector(0 downto 0);  -- Delay4:output -> cast182:input
	signal cast182_output_wire                      : std_logic;                     -- cast182:output -> Acc_Histogram:we
	signal counter_q_wire                           : std_logic_vector(19 downto 0); -- Counter:q -> cast183:input
	signal cast183_output_wire                      : std_logic_vector(20 downto 0); -- cast183:output -> Comparator:dataa
	signal cast184_output_wire                      : std_logic_vector(9 downto 0);  -- cast184:output -> Comparator1:dataa
	signal delay5_output_wire                       : std_logic_vector(9 downto 0);  -- Delay5:output -> cast185:input
	signal cast185_output_wire                      : std_logic_vector(7 downto 0);  -- cast185:output -> Acc_Histogram:write_address
	signal cast186_output_wire                      : std_logic_vector(10 downto 0); -- cast186:output -> Comparator6:dataa
	signal cast187_output_wire                      : std_logic_vector(10 downto 0); -- cast187:output -> Comparator7:dataa
	signal cast188_output_wire                      : std_logic_vector(10 downto 0); -- cast188:output -> Comparator8:dataa
	signal addr_in_0_output_wire                    : std_logic_vector(7 downto 0);  -- addr_in_0:output -> cast189:input
	signal cast189_output_wire                      : std_logic_vector(7 downto 0);  -- cast189:output -> Acc_Histogram:read_address
	signal cast190_output_wire                      : std_logic;                     -- cast190:output -> Counter2:cnt_ena
	signal cast191_output_wire                      : std_logic_vector(10 downto 0); -- cast191:output -> Comparator4:datab
	signal cast192_output_wire                      : std_logic_vector(8 downto 0);  -- cast192:output -> Comparator2:datab
	signal cast193_output_wire                      : std_logic_vector(8 downto 0);  -- cast193:output -> Comparator5:datab
	signal cast194_output_wire                      : std_logic_vector(10 downto 0); -- cast194:output -> Comparator4:dataa
	signal cast195_output_wire                      : std_logic_vector(15 downto 0); -- cast195:output -> Histogram:data
	signal multiplexer5_result_wire                 : std_logic_vector(9 downto 0);  -- Multiplexer5:result -> cast196:input
	signal cast196_output_wire                      : std_logic_vector(7 downto 0);  -- cast196:output -> Histogram:write_address
	signal multiplexer_result_wire                  : std_logic_vector(8 downto 0);  -- Multiplexer:result -> cast197:input
	signal cast197_output_wire                      : std_logic_vector(7 downto 0);  -- cast197:output -> Histogram:read_address
	signal multiplexer6_result_wire                 : std_logic_vector(0 downto 0);  -- Multiplexer6:result -> cast198:input
	signal cast198_output_wire                      : std_logic;                     -- cast198:output -> Histogram:we
	signal logical_bit_operator1_result_wire        : std_logic;                     -- Logical_Bit_Operator1:result -> cast199:input
	signal cast199_output_wire                      : std_logic_vector(0 downto 0);  -- cast199:output -> Delay:input
	signal cast200_output_wire                      : std_logic;                     -- cast200:output -> Logical_Bit_Operator6:data0
	signal logical_bit_operator7_result_wire        : std_logic;                     -- Logical_Bit_Operator7:result -> cast201:input
	signal cast201_output_wire                      : std_logic_vector(0 downto 0);  -- cast201:output -> Delay2:input
	signal cast202_output_wire                      : std_logic_vector(8 downto 0);  -- cast202:output -> Comparator2:dataa
	signal logical_bit_operator8_result_wire        : std_logic;                     -- Logical_Bit_Operator8:result -> cast203:input
	signal cast203_output_wire                      : std_logic_vector(0 downto 0);  -- cast203:output -> Memory_Delay3:input
	signal memory_delay4_output_wire                : std_logic_vector(7 downto 0);  -- Memory_Delay4:output -> cast204:input
	signal cast204_output_wire                      : std_logic_vector(8 downto 0);  -- cast204:output -> Comparator5:dataa
	signal logical_bit_operator10_result_wire       : std_logic;                     -- Logical_Bit_Operator10:result -> cast205:input
	signal cast205_output_wire                      : std_logic_vector(0 downto 0);  -- cast205:output -> Memory_Delay6:input
	signal cast206_output_wire                      : std_logic_vector(0 downto 0);  -- cast206:output -> Memory_Delay7:input
	signal cast207_output_wire                      : std_logic;                     -- cast207:output -> Logical_Bit_Operator8:data2
	signal memory_delay8_output_wire                : std_logic_vector(0 downto 0);  -- Memory_Delay8:output -> cast208:input
	signal cast208_output_wire                      : std_logic;                     -- cast208:output -> Logical_Bit_Operator10:data2
	signal cast209_output_wire                      : std_logic_vector(0 downto 0);  -- cast209:output -> Multiplexer:sel
	signal cast210_output_wire                      : std_logic_vector(8 downto 0);  -- cast210:output -> Multiplexer:in0
	signal comparator1_result_wire                  : std_logic;                     -- Comparator1:result -> cast211:input
	signal cast211_output_wire                      : std_logic_vector(0 downto 0);  -- cast211:output -> Multiplexer1:sel
	signal cast212_output_wire                      : std_logic_vector(10 downto 0); -- cast212:output -> Multiplexer1:in0
	signal comparator3_result_wire                  : std_logic;                     -- Comparator3:result -> cast213:input
	signal cast213_output_wire                      : std_logic_vector(0 downto 0);  -- cast213:output -> Multiplexer2:sel
	signal constant8_output_wire                    : std_logic_vector(7 downto 0);  -- Constant8:output -> cast214:input
	signal cast214_output_wire                      : std_logic_vector(10 downto 0); -- cast214:output -> Multiplexer2:in1
	signal constant9_output_wire                    : std_logic_vector(31 downto 0); -- Constant9:output -> cast215:input
	signal cast215_output_wire                      : std_logic_vector(55 downto 0); -- cast215:output -> Multiplexer3:in1
	signal cast216_output_wire                      : std_logic_vector(0 downto 0);  -- cast216:output -> Multiplexer4:sel
	signal cast217_output_wire                      : std_logic_vector(0 downto 0);  -- cast217:output -> Multiplexer5:sel
	signal memory_delay1_output_wire                : std_logic_vector(7 downto 0);  -- Memory_Delay1:output -> cast218:input
	signal cast218_output_wire                      : std_logic_vector(9 downto 0);  -- cast218:output -> Multiplexer5:in0
	signal cast219_output_wire                      : std_logic_vector(0 downto 0);  -- cast219:output -> Multiplexer6:sel
	signal cast220_output_wire                      : std_logic_vector(16 downto 0); -- cast220:output -> Multiplexer7:in1
	signal histogram_q_wire                         : std_logic_vector(15 downto 0); -- Histogram:q -> [cast221:input, cast223:input]
	signal cast221_output_wire                      : std_logic_vector(16 downto 0); -- cast221:output -> Multiplexer8:in0
	signal memory_delay5_output_wire                : std_logic_vector(15 downto 0); -- Memory_Delay5:output -> cast222:input
	signal cast222_output_wire                      : std_logic_vector(16 downto 0); -- cast222:output -> Multiplexer8:in1
	signal cast223_output_wire                      : std_logic_vector(15 downto 0); -- cast223:output -> Multiplier1:dataa
	signal multiplexer2_result_wire                 : std_logic_vector(10 downto 0); -- Multiplexer2:result -> [cast224:input, cast230:input]
	signal cast224_output_wire                      : std_logic_vector(7 downto 0);  -- cast224:output -> Multiplier1:datab
	signal multiplexer7_result_wire                 : std_logic_vector(16 downto 0); -- Multiplexer7:result -> cast225:input
	signal cast225_output_wire                      : std_logic_vector(15 downto 0); -- cast225:output -> Pipelined_Adder:dataa
	signal multiplier1_result_wire                  : std_logic_vector(23 downto 0); -- Multiplier1:result -> cast226:input
	signal cast226_output_wire                      : std_logic_vector(31 downto 0); -- cast226:output -> Pipelined_Adder1:dataa
	signal multiplexer3_result_wire                 : std_logic_vector(55 downto 0); -- Multiplexer3:result -> cast227:input
	signal cast227_output_wire                      : std_logic_vector(31 downto 0); -- cast227:output -> Pipelined_Adder1:datab
	signal pipelined_adder1_result_wire             : std_logic_vector(31 downto 0); -- Pipelined_Adder1:result -> [cast228:input, cast229:input]
	signal cast228_output_wire                      : std_logic_vector(31 downto 0); -- cast228:output -> Multiplier:dataa
	signal cast229_output_wire                      : std_logic_vector(55 downto 0); -- cast229:output -> Multiplexer3:in0
	signal cast230_output_wire                      : std_logic_vector(9 downto 0);  -- cast230:output -> Pipelined_Adder2:dataa
	signal pipelined_adder2_result_wire             : std_logic_vector(9 downto 0);  -- Pipelined_Adder2:result -> cast231:input
	signal cast231_output_wire                      : std_logic_vector(10 downto 0); -- cast231:output -> Multiplexer1:in1
	signal vcc_output_wire                          : std_logic;                     -- VCC:output -> cast232:input
	signal cast232_output_wire                      : std_logic_vector(0 downto 0);  -- cast232:output -> Multiplexer6:in1
	signal clock_0_clock_output_clk                 : std_logic;                     -- Clock_0:clock_out -> [Acc_Histogram:clock, Comparator1:clock, Comparator2:clock, Comparator3:clock, Comparator4:clock, Comparator5:clock, Comparator6:clock, Comparator7:clock, Comparator8:clock, Comparator:clock, Counter1:clock, Counter2:clock, Counter3:clock, Counter:clock, Delay1:clock, Delay2:clock, Delay4:clock, Delay5:clock, Delay:clock, Histogram:clock, Memory_Delay1:clock, Memory_Delay2:clock, Memory_Delay3:clock, Memory_Delay4:clock, Memory_Delay5:clock, Memory_Delay6:clock, Memory_Delay7:clock, Memory_Delay8:clock, Multiplexer1:clock, Multiplexer2:clock, Multiplexer3:clock, Multiplexer4:clock, Multiplexer5:clock, Multiplexer6:clock, Multiplexer7:clock, Multiplexer8:clock, Multiplexer:clock, Multiplier1:clock, Multiplier:clock, Pipelined_Adder1:clock, Pipelined_Adder2:clock, Pipelined_Adder:clock]
	signal clock_0_clock_output_reset               : std_logic;                     -- Clock_0:aclr_out -> [Comparator1:sclr, Comparator2:sclr, Comparator3:sclr, Comparator4:sclr, Comparator5:sclr, Comparator6:sclr, Comparator7:sclr, Comparator8:sclr, Comparator:sclr, Counter1:aclr, Counter2:aclr, Counter3:aclr, Counter:aclr, Delay1:aclr, Delay2:aclr, Delay4:aclr, Delay5:aclr, Delay:aclr, Memory_Delay1:aclr, Memory_Delay2:aclr, Memory_Delay3:aclr, Memory_Delay4:aclr, Memory_Delay5:aclr, Memory_Delay6:aclr, Memory_Delay7:aclr, Memory_Delay8:aclr, Multiplexer1:aclr, Multiplexer2:aclr, Multiplexer3:aclr, Multiplexer4:aclr, Multiplexer5:aclr, Multiplexer6:aclr, Multiplexer7:aclr, Multiplexer8:aclr, Multiplexer:aclr, Multiplier1:aclr, Multiplier:aclr, Pipelined_Adder1:aclr, Pipelined_Adder2:aclr, Pipelined_Adder:aclr]

begin

	clock_0 : component alt_dspbuilder_clock_GNQFU4PUDH
		port map (
			clock_out => clock_0_clock_output_clk,   -- clock_output.clk
			aclr_out  => clock_0_clock_output_reset, --             .reset
			clock     => Clock,                      --        clock.clk
			aclr      => reset                       --             .reset
		);

	valid_in_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => valid_in,               --  input.wire
			output => valid_in_0_output_wire  -- output.wire
		);

	multiplier1 : component alt_dspbuilder_multiplier_GNUSAT2VBO
		generic map (
			aWidth                         => 16,
			Signed                         => 0,
			bWidth                         => 8,
			DEDICATED_MULTIPLIER_CIRCUITRY => "YES",
			pipeline                       => 1,
			OutputLsb                      => 0,
			OutputMsb                      => 23
		)
		port map (
			clock     => clock_0_clock_output_clk,            -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,          --           .reset
			dataa     => cast223_output_wire,                 --      dataa.wire
			datab     => cast224_output_wire,                 --      datab.wire
			result    => multiplier1_result_wire,             --     result.wire
			user_aclr => multiplier1user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => multiplier1enavcc_output_wire        --        ena.wire
		);

	multiplier1user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplier1user_aclrgnd_output_wire  -- output.wire
		);

	multiplier1enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => multiplier1enavcc_output_wire  -- output.wire
		);

	binary_point_casting1 : component alt_dspbuilder_cast_GNBBMDRQ7A
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => cast175_output_wire,               --  input.wire
			output => binary_point_casting1_output_wire  -- output.wire
		);

	histogram : component dual_port_ram_sync
		port map (
			clock         => clock_0_clock_output_clk, --         clock.clk
			data          => cast195_output_wire,      --          data.wire
			write_address => cast196_output_wire,      -- write_address.wire
			read_address  => cast197_output_wire,      --  read_address.wire
			we            => cast198_output_wire,      --            we.wire
			q             => histogram_q_wire          --             q.wire
		);

	binary_point_casting2 : component alt_dspbuilder_cast_GNBBMDRQ7A
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => cast176_output_wire,               --  input.wire
			output => binary_point_casting2_output_wire  -- output.wire
		);

	multiplexer : component alt_dspbuilder_multiplexer_GNIM5IEXF4
		generic map (
			number_inputs          => 2,
			pipeline               => 0,
			width                  => 9,
			HDLTYPE                => "STD_LOGIC_VECTOR",
			use_one_hot_select_bus => 0
		)
		port map (
			clock     => clock_0_clock_output_clk,            -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,          --           .reset
			sel       => cast209_output_wire,                 --        sel.wire
			result    => multiplexer_result_wire,             --     result.wire
			ena       => multiplexerenavcc_output_wire,       --        ena.wire
			user_aclr => multiplexeruser_aclrgnd_output_wire, --  user_aclr.wire
			in0       => cast210_output_wire,                 --        in0.wire
			in1       => counter1_q_wire                      --        in1.wire
		);

	multiplexeruser_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplexeruser_aclrgnd_output_wire  -- output.wire
		);

	multiplexerenavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => multiplexerenavcc_output_wire  -- output.wire
		);

	pixel_in_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => pixel_in,               --  input.wire
			output => pixel_in_0_output_wire  -- output.wire
		);

	acc_histogram : component dual_port_ram_sync2
		port map (
			clock         => clock_0_clock_output_clk, --         clock.clk
			data          => cast174_output_wire,      --          data.wire
			write_address => cast185_output_wire,      -- write_address.wire
			read_address  => cast189_output_wire,      --  read_address.wire
			we            => cast182_output_wire,      --            we.wire
			q             => acc_histogram_q_wire,     --             q.wire
			max           => acc_histogram_max_wire    --           max.wire
		);

	delay : component alt_dspbuilder_delay_GNTBDM57LR
		generic map (
			ClockPhase => "1",
			BitPattern => "1",
			width      => 1,
			use_init   => 0,
			delay      => 2
		)
		port map (
			input  => cast199_output_wire,        --      input.wire
			clock  => clock_0_clock_output_clk,   -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset, --           .reset
			output => delay_output_wire,          --     output.wire
			sclr   => delaysclrgnd_output_wire,   --       sclr.wire
			ena    => delayenavcc_output_wire     --        ena.wire
		);

	delaysclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delaysclrgnd_output_wire  -- output.wire
		);

	delayenavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => delayenavcc_output_wire  -- output.wire
		);

	comparator : component alt_dspbuilder_comparator_GN
		generic map (
			Operator  => "Altagb",
			lpm_width => 21
		)
		port map (
			clock  => clock_0_clock_output_clk,   -- clock_sclr.clk
			sclr   => clock_0_clock_output_reset, --           .reset
			dataa  => cast183_output_wire,        --      dataa.wire
			datab  => cast177_output_wire,        --      datab.wire
			result => comparator_result_wire      --     result.wire
		);

	counter : component alt_dspbuilder_counter_GNS5ZU7DCJ
		generic map (
			svalue       => "1",
			use_cnt_ena  => "true",
			use_cout     => "false",
			modulus      => -1,
			use_sclr     => "true",
			ndirection   => 1,
			use_usr_aclr => "false",
			width        => 20,
			use_ena      => "false",
			use_sset     => "false",
			use_aload    => "false",
			avalue       => "0",
			use_aset     => "false",
			use_sload    => "false",
			use_cin      => "false"
		)
		port map (
			clock   => clock_0_clock_output_clk,          -- clock_aclr.clk
			aclr    => clock_0_clock_output_reset,        --           .reset
			cnt_ena => valid_in_0_output_wire,            --    cnt_ena.wire
			sclr    => logical_bit_operator5_result_wire, --       sclr.wire
			q       => counter_q_wire,                    --          q.wire
			cout    => open                               --       cout.wire
		);

	pipelined_adder2 : component alt_dspbuilder_pipelined_adder_GNY2JEH574
		generic map (
			pipeline => 0,
			width    => 10
		)
		port map (
			clock     => clock_0_clock_output_clk,                 -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,               --           .reset
			dataa     => cast230_output_wire,                      --      dataa.wire
			datab     => constant3_output_wire,                    --      datab.wire
			result    => pipelined_adder2_result_wire,             --     result.wire
			user_aclr => pipelined_adder2user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => pipelined_adder2enavcc_output_wire        --        ena.wire
		);

	pipelined_adder2user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => pipelined_adder2user_aclrgnd_output_wire  -- output.wire
		);

	pipelined_adder2enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => pipelined_adder2enavcc_output_wire  -- output.wire
		);

	pipelined_adder1 : component alt_dspbuilder_pipelined_adder_GNTWZRTG4I
		generic map (
			pipeline => 1,
			width    => 32
		)
		port map (
			clock     => clock_0_clock_output_clk,                 -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,               --           .reset
			dataa     => cast226_output_wire,                      --      dataa.wire
			datab     => cast227_output_wire,                      --      datab.wire
			result    => pipelined_adder1_result_wire,             --     result.wire
			user_aclr => pipelined_adder1user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => pipelined_adder1enavcc_output_wire        --        ena.wire
		);

	pipelined_adder1user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => pipelined_adder1user_aclrgnd_output_wire  -- output.wire
		);

	pipelined_adder1enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => pipelined_adder1enavcc_output_wire  -- output.wire
		);

	addr_in_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => addr_in,               --  input.wire
			output => addr_in_0_output_wire  -- output.wire
		);

	logical_bit_operator1 : component alt_dspbuilder_logical_bit_op_GNA5ZFEL7V
		generic map (
			LogicalOp     => "AltAND",
			number_inputs => 2
		)
		port map (
			result => logical_bit_operator1_result_wire, -- result.wire
			data0  => valid_in_0_output_wire,            --  data0.wire
			data1  => logical_bit_operator_result_wire   --  data1.wire
		);

	logical_bit_operator2 : component alt_dspbuilder_logical_bit_op_GNA5ZFEL7V
		generic map (
			LogicalOp     => "AltAND",
			number_inputs => 2
		)
		port map (
			result => logical_bit_operator2_result_wire, -- result.wire
			data0  => comparator_result_wire,            --  data0.wire
			data1  => comparator6_result_wire            --  data1.wire
		);

	max_out_0 : component alt_dspbuilder_port_GNEPKLLZKY
		port map (
			input  => binary_point_casting2_output_wire, --  input.wire
			output => max_out                            -- output.wire
		);

	logical_bit_operator3 : component alt_dspbuilder_logical_bit_op_GNA5ZFEL7V
		generic map (
			LogicalOp     => "AltAND",
			number_inputs => 2
		)
		port map (
			result => logical_bit_operator3_result_wire, -- result.wire
			data0  => comparator7_result_wire,           --  data0.wire
			data1  => comparator8_result_wire            --  data1.wire
		);

	constant2 : component alt_dspbuilder_constant_GNIIAAYRYZ
		generic map (
			BitPattern => "000000000000000000110110",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 24
		)
		port map (
			output => constant2_output_wire  -- output.wire
		);

	logical_bit_operator4 : component alt_dspbuilder_logical_bit_op_GNKUBZL4TE
		generic map (
			LogicalOp     => "AltNOT",
			number_inputs => 1
		)
		port map (
			result => logical_bit_operator4_result_wire, -- result.wire
			data0  => comparator8_result_wire            --  data0.wire
		);

	comparator8 : component alt_dspbuilder_comparator_GN
		generic map (
			Operator  => "Altalb",
			lpm_width => 11
		)
		port map (
			clock  => clock_0_clock_output_clk,   -- clock_sclr.clk
			sclr   => clock_0_clock_output_reset, --           .reset
			dataa  => cast188_output_wire,        --      dataa.wire
			datab  => cast180_output_wire,        --      datab.wire
			result => comparator8_result_wire     --     result.wire
		);

	constant3 : component alt_dspbuilder_constant_GNTHQFUUUC
		generic map (
			BitPattern => "0000000001",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 10
		)
		port map (
			output => constant3_output_wire  -- output.wire
		);

	logical_bit_operator5 : component alt_dspbuilder_logical_bit_op_GNA5ZFEL7V
		generic map (
			LogicalOp     => "AltAND",
			number_inputs => 2
		)
		port map (
			result => logical_bit_operator5_result_wire, -- result.wire
			data0  => eof_in_0_output_wire,              --  data0.wire
			data1  => logical_bit_operator4_result_wire  --  data1.wire
		);

	comparator7 : component alt_dspbuilder_comparator_GN
		generic map (
			Operator  => "Altagb",
			lpm_width => 11
		)
		port map (
			clock  => clock_0_clock_output_clk,   -- clock_sclr.clk
			sclr   => clock_0_clock_output_reset, --           .reset
			dataa  => cast187_output_wire,        --      dataa.wire
			datab  => cast179_output_wire,        --      datab.wire
			result => comparator7_result_wire     --     result.wire
		);

	logical_bit_operator6 : component alt_dspbuilder_logical_bit_op_GNUQ2R64DV
		generic map (
			LogicalOp     => "AltOR",
			number_inputs => 2
		)
		port map (
			result => logical_bit_operator6_result_wire, -- result.wire
			data0  => cast200_output_wire,               --  data0.wire
			data1  => logical_bit_operator5_result_wire  --  data1.wire
		);

	comparator6 : component alt_dspbuilder_comparator_GN
		generic map (
			Operator  => "Altalb",
			lpm_width => 11
		)
		port map (
			clock  => clock_0_clock_output_clk,   -- clock_sclr.clk
			sclr   => clock_0_clock_output_reset, --           .reset
			dataa  => cast186_output_wire,        --      dataa.wire
			datab  => cast178_output_wire,        --      datab.wire
			result => comparator6_result_wire     --     result.wire
		);

	constant1 : component alt_dspbuilder_constant_GNLUER2G5H
		generic map (
			BitPattern => "1001010111111111111",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 19
		)
		port map (
			output => constant1_output_wire  -- output.wire
		);

	logical_bit_operator10 : component alt_dspbuilder_logical_bit_op_GN5A3KLAEC
		generic map (
			LogicalOp     => "AltAND",
			number_inputs => 3
		)
		port map (
			result => logical_bit_operator10_result_wire, -- result.wire
			data0  => comparator5_result_wire,            --  data0.wire
			data1  => valid_in_0_output_wire,             --  data1.wire
			data2  => cast208_output_wire                 --  data2.wire
		);

	logical_bit_operator7 : component alt_dspbuilder_logical_bit_op_GNA5ZFEL7V
		generic map (
			LogicalOp     => "AltAND",
			number_inputs => 2
		)
		port map (
			result => logical_bit_operator7_result_wire, -- result.wire
			data0  => comparator_result_wire,            --  data0.wire
			data1  => comparator4_result_wire            --  data1.wire
		);

	logical_bit_operator8 : component alt_dspbuilder_logical_bit_op_GN5A3KLAEC
		generic map (
			LogicalOp     => "AltAND",
			number_inputs => 3
		)
		port map (
			result => logical_bit_operator8_result_wire, -- result.wire
			data0  => comparator2_result_wire,           --  data0.wire
			data1  => valid_in_0_output_wire,            --  data1.wire
			data2  => cast207_output_wire                --  data2.wire
		);

	constant8 : component alt_dspbuilder_constant_GNC5NOVIJT
		generic map (
			BitPattern => "00000000",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 8
		)
		port map (
			output => constant8_output_wire  -- output.wire
		);

	constant9 : component alt_dspbuilder_constant_GNRSDUIWRP
		generic map (
			BitPattern => "00000000000000000000000000000000",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 32
		)
		port map (
			output => constant9_output_wire  -- output.wire
		);

	constant7 : component alt_dspbuilder_constant_GN5IRMZXKK
		generic map (
			BitPattern => "0000000000",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 10
		)
		port map (
			output => constant7_output_wire  -- output.wire
		);

	constant4 : component alt_dspbuilder_constant_GNWFCSDEFM
		generic map (
			BitPattern => "0000000000000001",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 16
		)
		port map (
			output => constant4_output_wire  -- output.wire
		);

	constant5 : component alt_dspbuilder_constant_GN5IRMZXKK
		generic map (
			BitPattern => "0000000000",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 10
		)
		port map (
			output => constant5_output_wire  -- output.wire
		);

	vcc : component alt_dspbuilder_vcc_GN
		port map (
			output => vcc_output_wire  -- output.wire
		);

	logical_bit_operator : component alt_dspbuilder_logical_bit_op_GNKUBZL4TE
		generic map (
			LogicalOp     => "AltNOT",
			number_inputs => 1
		)
		port map (
			result => logical_bit_operator_result_wire, -- result.wire
			data0  => comparator_result_wire            --  data0.wire
		);

	multiplexer3 : component alt_dspbuilder_multiplexer_GNTG7F5PN7
		generic map (
			number_inputs          => 2,
			pipeline               => 0,
			width                  => 56,
			HDLTYPE                => "STD_LOGIC_VECTOR",
			use_one_hot_select_bus => 0
		)
		port map (
			clock     => clock_0_clock_output_clk,             -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,           --           .reset
			sel       => delay1_output_wire,                   --        sel.wire
			result    => multiplexer3_result_wire,             --     result.wire
			ena       => multiplexer3enavcc_output_wire,       --        ena.wire
			user_aclr => multiplexer3user_aclrgnd_output_wire, --  user_aclr.wire
			in0       => cast229_output_wire,                  --        in0.wire
			in1       => cast215_output_wire                   --        in1.wire
		);

	multiplexer3user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplexer3user_aclrgnd_output_wire  -- output.wire
		);

	multiplexer3enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => multiplexer3enavcc_output_wire  -- output.wire
		);

	multiplexer4 : component alt_dspbuilder_multiplexer_GN7X7SG76C
		generic map (
			number_inputs          => 2,
			pipeline               => 0,
			width                  => 16,
			HDLTYPE                => "STD_LOGIC_VECTOR",
			use_one_hot_select_bus => 0
		)
		port map (
			clock     => clock_0_clock_output_clk,             -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,           --           .reset
			sel       => cast216_output_wire,                  --        sel.wire
			result    => multiplexer4_result_wire,             --     result.wire
			ena       => multiplexer4enavcc_output_wire,       --        ena.wire
			user_aclr => multiplexer4user_aclrgnd_output_wire, --  user_aclr.wire
			in0       => pipelined_adder_result_wire,          --        in0.wire
			in1       => constant13_output_wire                --        in1.wire
		);

	multiplexer4user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplexer4user_aclrgnd_output_wire  -- output.wire
		);

	multiplexer4enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => multiplexer4enavcc_output_wire  -- output.wire
		);

	multiplexer1 : component alt_dspbuilder_multiplexer_GNCMV7Z7A7
		generic map (
			number_inputs          => 2,
			pipeline               => 1,
			width                  => 11,
			HDLTYPE                => "STD_LOGIC_VECTOR",
			use_one_hot_select_bus => 0
		)
		port map (
			clock     => clock_0_clock_output_clk,             -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,           --           .reset
			sel       => cast211_output_wire,                  --        sel.wire
			result    => multiplexer1_result_wire,             --     result.wire
			ena       => multiplexer1enavcc_output_wire,       --        ena.wire
			user_aclr => multiplexer1user_aclrgnd_output_wire, --  user_aclr.wire
			in0       => cast212_output_wire,                  --        in0.wire
			in1       => cast231_output_wire                   --        in1.wire
		);

	multiplexer1user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplexer1user_aclrgnd_output_wire  -- output.wire
		);

	multiplexer1enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => multiplexer1enavcc_output_wire  -- output.wire
		);

	multiplexer2 : component alt_dspbuilder_multiplexer_GNXY3BAFE2
		generic map (
			number_inputs          => 2,
			pipeline               => 0,
			width                  => 11,
			HDLTYPE                => "STD_LOGIC_VECTOR",
			use_one_hot_select_bus => 0
		)
		port map (
			clock     => clock_0_clock_output_clk,             -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,           --           .reset
			sel       => cast213_output_wire,                  --        sel.wire
			result    => multiplexer2_result_wire,             --     result.wire
			ena       => multiplexer2enavcc_output_wire,       --        ena.wire
			user_aclr => multiplexer2user_aclrgnd_output_wire, --  user_aclr.wire
			in0       => multiplexer1_result_wire,             --        in0.wire
			in1       => cast214_output_wire                   --        in1.wire
		);

	multiplexer2user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplexer2user_aclrgnd_output_wire  -- output.wire
		);

	multiplexer2enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => multiplexer2enavcc_output_wire  -- output.wire
		);

	memory_delay7 : component alt_dspbuilder_memdelay_GNSNJI6FHR
		generic map (
			RAMTYPE => "AUTO",
			WIDTH   => 1,
			DELAY   => 1
		)
		port map (
			clock     => clock_0_clock_output_clk,              -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,            --           .reset
			input     => cast206_output_wire,                   --      input.wire
			output    => memory_delay7_output_wire,             --     output.wire
			user_aclr => memory_delay7user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => memory_delay7enavcc_output_wire        --        ena.wire
		);

	memory_delay7user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => memory_delay7user_aclrgnd_output_wire  -- output.wire
		);

	memory_delay7enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => memory_delay7enavcc_output_wire  -- output.wire
		);

	pipelined_adder : component alt_dspbuilder_pipelined_adder_GNTWZRTG4I
		generic map (
			pipeline => 1,
			width    => 16
		)
		port map (
			clock     => clock_0_clock_output_clk,                -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,              --           .reset
			dataa     => cast225_output_wire,                     --      dataa.wire
			datab     => constant4_output_wire,                   --      datab.wire
			result    => pipelined_adder_result_wire,             --     result.wire
			user_aclr => pipelined_adderuser_aclrgnd_output_wire, --  user_aclr.wire
			ena       => pipelined_adderenavcc_output_wire        --        ena.wire
		);

	pipelined_adderuser_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => pipelined_adderuser_aclrgnd_output_wire  -- output.wire
		);

	pipelined_adderenavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => pipelined_adderenavcc_output_wire  -- output.wire
		);

	memory_delay8 : component alt_dspbuilder_memdelay_GNSNJI6FHR
		generic map (
			RAMTYPE => "AUTO",
			WIDTH   => 1,
			DELAY   => 1
		)
		port map (
			clock     => clock_0_clock_output_clk,              -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,            --           .reset
			input     => memory_delay7_output_wire,             --      input.wire
			output    => memory_delay8_output_wire,             --     output.wire
			user_aclr => memory_delay8user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => memory_delay8enavcc_output_wire        --        ena.wire
		);

	memory_delay8user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => memory_delay8user_aclrgnd_output_wire  -- output.wire
		);

	memory_delay8enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => memory_delay8enavcc_output_wire  -- output.wire
		);

	memory_delay5 : component alt_dspbuilder_memdelay_GNMIZKWFE6
		generic map (
			RAMTYPE => "AUTO",
			WIDTH   => 16,
			DELAY   => 1
		)
		port map (
			clock     => clock_0_clock_output_clk,              -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,            --           .reset
			input     => multiplexer4_result_wire,              --      input.wire
			output    => memory_delay5_output_wire,             --     output.wire
			user_aclr => memory_delay5user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => memory_delay5enavcc_output_wire        --        ena.wire
		);

	memory_delay5user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => memory_delay5user_aclrgnd_output_wire  -- output.wire
		);

	memory_delay5enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => memory_delay5enavcc_output_wire  -- output.wire
		);

	memory_delay6 : component alt_dspbuilder_memdelay_GNSNJI6FHR
		generic map (
			RAMTYPE => "AUTO",
			WIDTH   => 1,
			DELAY   => 1
		)
		port map (
			clock     => clock_0_clock_output_clk,              -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,            --           .reset
			input     => cast205_output_wire,                   --      input.wire
			output    => memory_delay6_output_wire,             --     output.wire
			user_aclr => memory_delay6user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => memory_delay6enavcc_output_wire        --        ena.wire
		);

	memory_delay6user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => memory_delay6user_aclrgnd_output_wire  -- output.wire
		);

	memory_delay6enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => memory_delay6enavcc_output_wire  -- output.wire
		);

	comparator1 : component alt_dspbuilder_comparator_GN
		generic map (
			Operator  => "Altagb",
			lpm_width => 10
		)
		port map (
			clock  => clock_0_clock_output_clk,   -- clock_sclr.clk
			sclr   => clock_0_clock_output_reset, --           .reset
			dataa  => cast184_output_wire,        --      dataa.wire
			datab  => constant5_output_wire,      --      datab.wire
			result => comparator1_result_wire     --     result.wire
		);

	comparator5 : component alt_dspbuilder_comparator_GN
		generic map (
			Operator  => "Altaeb",
			lpm_width => 9
		)
		port map (
			clock  => clock_0_clock_output_clk,   -- clock_sclr.clk
			sclr   => clock_0_clock_output_reset, --           .reset
			dataa  => cast204_output_wire,        --      dataa.wire
			datab  => cast193_output_wire,        --      datab.wire
			result => comparator5_result_wire     --     result.wire
		);

	memory_delay3 : component alt_dspbuilder_memdelay_GNSNJI6FHR
		generic map (
			RAMTYPE => "AUTO",
			WIDTH   => 1,
			DELAY   => 1
		)
		port map (
			clock     => clock_0_clock_output_clk,              -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,            --           .reset
			input     => cast203_output_wire,                   --      input.wire
			output    => memory_delay3_output_wire,             --     output.wire
			user_aclr => memory_delay3user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => memory_delay3enavcc_output_wire        --        ena.wire
		);

	memory_delay3user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => memory_delay3user_aclrgnd_output_wire  -- output.wire
		);

	memory_delay3enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => memory_delay3enavcc_output_wire  -- output.wire
		);

	comparator4 : component alt_dspbuilder_comparator_GN
		generic map (
			Operator  => "Altaeb",
			lpm_width => 11
		)
		port map (
			clock  => clock_0_clock_output_clk,   -- clock_sclr.clk
			sclr   => clock_0_clock_output_reset, --           .reset
			dataa  => cast194_output_wire,        --      dataa.wire
			datab  => cast191_output_wire,        --      datab.wire
			result => comparator4_result_wire     --     result.wire
		);

	memory_delay4 : component alt_dspbuilder_memdelay_GN7KC3ZSDB
		generic map (
			RAMTYPE => "AUTO",
			WIDTH   => 8,
			DELAY   => 1
		)
		port map (
			clock     => clock_0_clock_output_clk,              -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,            --           .reset
			input     => memory_delay2_output_wire,             --      input.wire
			output    => memory_delay4_output_wire,             --     output.wire
			user_aclr => memory_delay4user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => memory_delay4enavcc_output_wire        --        ena.wire
		);

	memory_delay4user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => memory_delay4user_aclrgnd_output_wire  -- output.wire
		);

	memory_delay4enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => memory_delay4enavcc_output_wire  -- output.wire
		);

	comparator3 : component alt_dspbuilder_comparator_GN
		generic map (
			Operator  => "Altalb",
			lpm_width => 11
		)
		port map (
			clock  => clock_0_clock_output_clk,   -- clock_sclr.clk
			sclr   => clock_0_clock_output_reset, --           .reset
			dataa  => multiplexer1_result_wire,   --      dataa.wire
			datab  => cast181_output_wire,        --      datab.wire
			result => comparator3_result_wire     --     result.wire
		);

	memory_delay1 : component alt_dspbuilder_memdelay_GNXMJOJMJV
		generic map (
			RAMTYPE => "AUTO",
			WIDTH   => 8,
			DELAY   => 2
		)
		port map (
			clock     => clock_0_clock_output_clk,              -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,            --           .reset
			input     => pixel_in_0_output_wire,                --      input.wire
			output    => memory_delay1_output_wire,             --     output.wire
			user_aclr => memory_delay1user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => memory_delay1enavcc_output_wire        --        ena.wire
		);

	memory_delay1user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => memory_delay1user_aclrgnd_output_wire  -- output.wire
		);

	memory_delay1enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => memory_delay1enavcc_output_wire  -- output.wire
		);

	comparator2 : component alt_dspbuilder_comparator_GN
		generic map (
			Operator  => "Altaeb",
			lpm_width => 9
		)
		port map (
			clock  => clock_0_clock_output_clk,   -- clock_sclr.clk
			sclr   => clock_0_clock_output_reset, --           .reset
			dataa  => cast202_output_wire,        --      dataa.wire
			datab  => cast192_output_wire,        --      datab.wire
			result => comparator2_result_wire     --     result.wire
		);

	memory_delay2 : component alt_dspbuilder_memdelay_GN7KC3ZSDB
		generic map (
			RAMTYPE => "AUTO",
			WIDTH   => 8,
			DELAY   => 1
		)
		port map (
			clock     => clock_0_clock_output_clk,              -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,            --           .reset
			input     => pixel_in_0_output_wire,                --      input.wire
			output    => memory_delay2_output_wire,             --     output.wire
			user_aclr => memory_delay2user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => memory_delay2enavcc_output_wire        --        ena.wire
		);

	memory_delay2user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => memory_delay2user_aclrgnd_output_wire  -- output.wire
		);

	memory_delay2enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => memory_delay2enavcc_output_wire  -- output.wire
		);

	multiplier : component alt_dspbuilder_multiplier_GNXX7E2RLJ
		generic map (
			aWidth                         => 32,
			Signed                         => 0,
			bWidth                         => 24,
			DEDICATED_MULTIPLIER_CIRCUITRY => "YES",
			pipeline                       => 1,
			OutputLsb                      => 0,
			OutputMsb                      => 31
		)
		port map (
			clock     => clock_0_clock_output_clk,           -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,         --           .reset
			dataa     => cast228_output_wire,                --      dataa.wire
			datab     => constant2_output_wire,              --      datab.wire
			result    => multiplier_result_wire,             --     result.wire
			user_aclr => multiplieruser_aclrgnd_output_wire, --  user_aclr.wire
			ena       => multiplierenavcc_output_wire        --        ena.wire
		);

	multiplieruser_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplieruser_aclrgnd_output_wire  -- output.wire
		);

	multiplierenavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => multiplierenavcc_output_wire  -- output.wire
		);

	value_out_0 : component alt_dspbuilder_port_GNEPKLLZKY
		port map (
			input  => binary_point_casting1_output_wire, --  input.wire
			output => value_out                          -- output.wire
		);

	delay2 : component alt_dspbuilder_delay_GNGQ56ZS4N
		generic map (
			ClockPhase => "1",
			BitPattern => "1",
			width      => 1,
			use_init   => 0,
			delay      => 1
		)
		port map (
			input  => cast201_output_wire,        --      input.wire
			clock  => clock_0_clock_output_clk,   -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset, --           .reset
			output => delay2_output_wire,         --     output.wire
			sclr   => delay2sclrgnd_output_wire,  --       sclr.wire
			ena    => delay2enavcc_output_wire    --        ena.wire
		);

	delay2sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delay2sclrgnd_output_wire  -- output.wire
		);

	delay2enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => delay2enavcc_output_wire  -- output.wire
		);

	delay1 : component alt_dspbuilder_delay_GNNQSQIG3K
		generic map (
			ClockPhase => "1",
			BitPattern => "1",
			width      => 1,
			use_init   => 0,
			delay      => 3
		)
		port map (
			input  => delay2_output_wire,         --      input.wire
			clock  => clock_0_clock_output_clk,   -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset, --           .reset
			output => delay1_output_wire,         --     output.wire
			sclr   => delay1sclrgnd_output_wire,  --       sclr.wire
			ena    => delay1enavcc_output_wire    --        ena.wire
		);

	delay1sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delay1sclrgnd_output_wire  -- output.wire
		);

	delay1enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => delay1enavcc_output_wire  -- output.wire
		);

	constant14 : component alt_dspbuilder_constant_GNQE5XU76S
		generic map (
			BitPattern => "0100000000",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 10
		)
		port map (
			output => constant14_output_wire  -- output.wire
		);

	constant13 : component alt_dspbuilder_constant_GNCWI5QDAD
		generic map (
			BitPattern => "0000000000000000",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 16
		)
		port map (
			output => constant13_output_wire  -- output.wire
		);

	constant12 : component alt_dspbuilder_constant_GNK57PM5EK
		generic map (
			BitPattern => "0011111111",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 10
		)
		port map (
			output => constant12_output_wire  -- output.wire
		);

	constant11 : component alt_dspbuilder_constant_GNSXLT2IGA
		generic map (
			BitPattern => "100000000",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 9
		)
		port map (
			output => constant11_output_wire  -- output.wire
		);

	eof_in_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => eof_in,               --  input.wire
			output => eof_in_0_output_wire  -- output.wire
		);

	binary_point_casting : component alt_dspbuilder_cast_GNBBMDRQ7A
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => multiplier_result_wire,           --  input.wire
			output => binary_point_casting_output_wire  -- output.wire
		);

	counter1 : component alt_dspbuilder_counter_GNJYRI37NB
		generic map (
			svalue       => "1",
			use_cnt_ena  => "true",
			use_cout     => "false",
			modulus      => -1,
			use_sclr     => "true",
			ndirection   => 1,
			use_usr_aclr => "false",
			width        => 9,
			use_ena      => "false",
			use_sset     => "false",
			use_aload    => "false",
			avalue       => "0",
			use_aset     => "false",
			use_sload    => "false",
			use_cin      => "false"
		)
		port map (
			clock   => clock_0_clock_output_clk,          -- clock_aclr.clk
			aclr    => clock_0_clock_output_reset,        --           .reset
			cnt_ena => logical_bit_operator2_result_wire, --    cnt_ena.wire
			sclr    => logical_bit_operator6_result_wire, --       sclr.wire
			q       => counter1_q_wire,                   --          q.wire
			cout    => open                               --       cout.wire
		);

	multiplexer7 : component alt_dspbuilder_multiplexer_GNMRY6PWYH
		generic map (
			number_inputs          => 2,
			pipeline               => 0,
			width                  => 17,
			HDLTYPE                => "STD_LOGIC_VECTOR",
			use_one_hot_select_bus => 0
		)
		port map (
			clock     => clock_0_clock_output_clk,             -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,           --           .reset
			sel       => memory_delay3_output_wire,            --        sel.wire
			result    => multiplexer7_result_wire,             --     result.wire
			ena       => multiplexer7enavcc_output_wire,       --        ena.wire
			user_aclr => multiplexer7user_aclrgnd_output_wire, --  user_aclr.wire
			in0       => multiplexer8_result_wire,             --        in0.wire
			in1       => cast220_output_wire                   --        in1.wire
		);

	multiplexer7user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplexer7user_aclrgnd_output_wire  -- output.wire
		);

	multiplexer7enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => multiplexer7enavcc_output_wire  -- output.wire
		);

	delay5 : component alt_dspbuilder_delay_GNUACQWN66
		generic map (
			ClockPhase => "1",
			BitPattern => "0000000001",
			width      => 10,
			use_init   => 0,
			delay      => 4
		)
		port map (
			input  => counter2_q_wire,            --      input.wire
			clock  => clock_0_clock_output_clk,   -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset, --           .reset
			output => delay5_output_wire,         --     output.wire
			sclr   => delay5sclrgnd_output_wire,  --       sclr.wire
			ena    => delay5enavcc_output_wire    --        ena.wire
		);

	delay5sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delay5sclrgnd_output_wire  -- output.wire
		);

	delay5enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => delay5enavcc_output_wire  -- output.wire
		);

	multiplexer8 : component alt_dspbuilder_multiplexer_GNMRY6PWYH
		generic map (
			number_inputs          => 2,
			pipeline               => 0,
			width                  => 17,
			HDLTYPE                => "STD_LOGIC_VECTOR",
			use_one_hot_select_bus => 0
		)
		port map (
			clock     => clock_0_clock_output_clk,             -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,           --           .reset
			sel       => memory_delay6_output_wire,            --        sel.wire
			result    => multiplexer8_result_wire,             --     result.wire
			ena       => multiplexer8enavcc_output_wire,       --        ena.wire
			user_aclr => multiplexer8user_aclrgnd_output_wire, --  user_aclr.wire
			in0       => cast221_output_wire,                  --        in0.wire
			in1       => cast222_output_wire                   --        in1.wire
		);

	multiplexer8user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplexer8user_aclrgnd_output_wire  -- output.wire
		);

	multiplexer8enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => multiplexer8enavcc_output_wire  -- output.wire
		);

	counter3 : component alt_dspbuilder_counter_GNPVW56BJJ
		generic map (
			svalue       => "1",
			use_cnt_ena  => "true",
			use_cout     => "false",
			modulus      => -1,
			use_sclr     => "true",
			ndirection   => 1,
			use_usr_aclr => "false",
			width        => 10,
			use_ena      => "false",
			use_sset     => "false",
			use_aload    => "false",
			avalue       => "0",
			use_aset     => "false",
			use_sload    => "false",
			use_cin      => "false"
		)
		port map (
			clock   => clock_0_clock_output_clk,          -- clock_aclr.clk
			aclr    => clock_0_clock_output_reset,        --           .reset
			cnt_ena => logical_bit_operator3_result_wire, --    cnt_ena.wire
			sclr    => logical_bit_operator5_result_wire, --       sclr.wire
			q       => counter3_q_wire,                   --          q.wire
			cout    => open                               --       cout.wire
		);

	delay4 : component alt_dspbuilder_delay_GNQBXYU75H
		generic map (
			ClockPhase => "1",
			BitPattern => "1",
			width      => 1,
			use_init   => 0,
			delay      => 4
		)
		port map (
			input  => delay2_output_wire,         --      input.wire
			clock  => clock_0_clock_output_clk,   -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset, --           .reset
			output => delay4_output_wire,         --     output.wire
			sclr   => delay4sclrgnd_output_wire,  --       sclr.wire
			ena    => delay4enavcc_output_wire    --        ena.wire
		);

	delay4sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delay4sclrgnd_output_wire  -- output.wire
		);

	delay4enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => delay4enavcc_output_wire  -- output.wire
		);

	multiplexer5 : component alt_dspbuilder_multiplexer_GNWZZP2IFI
		generic map (
			number_inputs          => 2,
			pipeline               => 0,
			width                  => 10,
			HDLTYPE                => "STD_LOGIC_VECTOR",
			use_one_hot_select_bus => 0
		)
		port map (
			clock     => clock_0_clock_output_clk,             -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,           --           .reset
			sel       => cast217_output_wire,                  --        sel.wire
			result    => multiplexer5_result_wire,             --     result.wire
			ena       => multiplexer5enavcc_output_wire,       --        ena.wire
			user_aclr => multiplexer5user_aclrgnd_output_wire, --  user_aclr.wire
			in0       => cast218_output_wire,                  --        in0.wire
			in1       => counter3_q_wire                       --        in1.wire
		);

	multiplexer5user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplexer5user_aclrgnd_output_wire  -- output.wire
		);

	multiplexer5enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => multiplexer5enavcc_output_wire  -- output.wire
		);

	counter2 : component alt_dspbuilder_counter_GNPVW56BJJ
		generic map (
			svalue       => "1",
			use_cnt_ena  => "true",
			use_cout     => "false",
			modulus      => -1,
			use_sclr     => "true",
			ndirection   => 1,
			use_usr_aclr => "false",
			width        => 10,
			use_ena      => "false",
			use_sset     => "false",
			use_aload    => "false",
			avalue       => "0",
			use_aset     => "false",
			use_sload    => "false",
			use_cin      => "false"
		)
		port map (
			clock   => clock_0_clock_output_clk,          -- clock_aclr.clk
			aclr    => clock_0_clock_output_reset,        --           .reset
			cnt_ena => cast190_output_wire,               --    cnt_ena.wire
			sclr    => logical_bit_operator5_result_wire, --       sclr.wire
			q       => counter2_q_wire,                   --          q.wire
			cout    => open                               --       cout.wire
		);

	multiplexer6 : component alt_dspbuilder_multiplexer_GNAIWAHV3K
		generic map (
			number_inputs          => 2,
			pipeline               => 0,
			width                  => 1,
			HDLTYPE                => "STD_LOGIC_VECTOR",
			use_one_hot_select_bus => 0
		)
		port map (
			clock     => clock_0_clock_output_clk,             -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,           --           .reset
			sel       => cast219_output_wire,                  --        sel.wire
			result    => multiplexer6_result_wire,             --     result.wire
			ena       => multiplexer6enavcc_output_wire,       --        ena.wire
			user_aclr => multiplexer6user_aclrgnd_output_wire, --  user_aclr.wire
			in0       => delay_output_wire,                    --        in0.wire
			in1       => cast232_output_wire                   --        in1.wire
		);

	multiplexer6user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplexer6user_aclrgnd_output_wire  -- output.wire
		);

	multiplexer6enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => multiplexer6enavcc_output_wire  -- output.wire
		);

	cast174 : component alt_dspbuilder_cast_GNU3FOKJ6W
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => binary_point_casting_output_wire, --  input.wire
			output => cast174_output_wire               -- output.wire
		);

	cast175 : component alt_dspbuilder_cast_GNHIWMUP5U
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => acc_histogram_q_wire, --  input.wire
			output => cast175_output_wire   -- output.wire
		);

	cast176 : component alt_dspbuilder_cast_GNHIWMUP5U
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => acc_histogram_max_wire, --  input.wire
			output => cast176_output_wire     -- output.wire
		);

	cast177 : component alt_dspbuilder_cast_GNOFO5NIX3
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => constant1_output_wire, --  input.wire
			output => cast177_output_wire    -- output.wire
		);

	cast178 : component alt_dspbuilder_cast_GN6OFM6A6B
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => constant11_output_wire, --  input.wire
			output => cast178_output_wire     -- output.wire
		);

	cast179 : component alt_dspbuilder_cast_GN5D52DF5S
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => constant12_output_wire, --  input.wire
			output => cast179_output_wire     -- output.wire
		);

	cast180 : component alt_dspbuilder_cast_GN5D52DF5S
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => constant14_output_wire, --  input.wire
			output => cast180_output_wire     -- output.wire
		);

	cast181 : component alt_dspbuilder_cast_GNAMS3PPNH
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => constant7_output_wire, --  input.wire
			output => cast181_output_wire    -- output.wire
		);

	cast182 : component alt_dspbuilder_cast_GNSB3OXIQS
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => delay4_output_wire,  --  input.wire
			output => cast182_output_wire  -- output.wire
		);

	cast183 : component alt_dspbuilder_cast_GN5JC4724B
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => counter_q_wire,      --  input.wire
			output => cast183_output_wire  -- output.wire
		);

	cast184 : component alt_dspbuilder_cast_GNPFJ7B3O7
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => counter1_q_wire,     --  input.wire
			output => cast184_output_wire  -- output.wire
		);

	cast185 : component alt_dspbuilder_cast_GNVKZTMEYW
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => delay5_output_wire,  --  input.wire
			output => cast185_output_wire  -- output.wire
		);

	cast186 : component alt_dspbuilder_cast_GN5D52DF5S
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => counter2_q_wire,     --  input.wire
			output => cast186_output_wire  -- output.wire
		);

	cast187 : component alt_dspbuilder_cast_GN5D52DF5S
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => counter2_q_wire,     --  input.wire
			output => cast187_output_wire  -- output.wire
		);

	cast188 : component alt_dspbuilder_cast_GN5D52DF5S
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => counter3_q_wire,     --  input.wire
			output => cast188_output_wire  -- output.wire
		);

	cast189 : component alt_dspbuilder_cast_GNBZR5PMEK
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => addr_in_0_output_wire, --  input.wire
			output => cast189_output_wire    -- output.wire
		);

	cast190 : component alt_dspbuilder_cast_GNSB3OXIQS
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => delay2_output_wire,  --  input.wire
			output => cast190_output_wire  -- output.wire
		);

	cast191 : component alt_dspbuilder_cast_GN5D52DF5S
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => counter2_q_wire,     --  input.wire
			output => cast191_output_wire  -- output.wire
		);

	cast192 : component alt_dspbuilder_cast_GNUW2C7J4Q
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => pixel_in_0_output_wire, --  input.wire
			output => cast192_output_wire     -- output.wire
		);

	cast193 : component alt_dspbuilder_cast_GNUW2C7J4Q
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => pixel_in_0_output_wire, --  input.wire
			output => cast193_output_wire     -- output.wire
		);

	cast194 : component alt_dspbuilder_cast_GN6OFM6A6B
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => counter1_q_wire,     --  input.wire
			output => cast194_output_wire  -- output.wire
		);

	cast195 : component alt_dspbuilder_cast_GNQQ42CR65
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => multiplexer4_result_wire, --  input.wire
			output => cast195_output_wire       -- output.wire
		);

	cast196 : component alt_dspbuilder_cast_GNVKZTMEYW
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => multiplexer5_result_wire, --  input.wire
			output => cast196_output_wire       -- output.wire
		);

	cast197 : component alt_dspbuilder_cast_GNSKTJRCBQ
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => multiplexer_result_wire, --  input.wire
			output => cast197_output_wire      -- output.wire
		);

	cast198 : component alt_dspbuilder_cast_GNSB3OXIQS
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => multiplexer6_result_wire, --  input.wire
			output => cast198_output_wire       -- output.wire
		);

	cast199 : component alt_dspbuilder_cast_GN46N4UJ5S
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => logical_bit_operator1_result_wire, --  input.wire
			output => cast199_output_wire                -- output.wire
		);

	cast200 : component alt_dspbuilder_cast_GNSB3OXIQS
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => delay2_output_wire,  --  input.wire
			output => cast200_output_wire  -- output.wire
		);

	cast201 : component alt_dspbuilder_cast_GN46N4UJ5S
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => logical_bit_operator7_result_wire, --  input.wire
			output => cast201_output_wire                -- output.wire
		);

	cast202 : component alt_dspbuilder_cast_GNUW2C7J4Q
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => memory_delay2_output_wire, --  input.wire
			output => cast202_output_wire        -- output.wire
		);

	cast203 : component alt_dspbuilder_cast_GN46N4UJ5S
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => logical_bit_operator8_result_wire, --  input.wire
			output => cast203_output_wire                -- output.wire
		);

	cast204 : component alt_dspbuilder_cast_GNUW2C7J4Q
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => memory_delay4_output_wire, --  input.wire
			output => cast204_output_wire        -- output.wire
		);

	cast205 : component alt_dspbuilder_cast_GN46N4UJ5S
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => logical_bit_operator10_result_wire, --  input.wire
			output => cast205_output_wire                 -- output.wire
		);

	cast206 : component alt_dspbuilder_cast_GN46N4UJ5S
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => valid_in_0_output_wire, --  input.wire
			output => cast206_output_wire     -- output.wire
		);

	cast207 : component alt_dspbuilder_cast_GNSB3OXIQS
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => memory_delay7_output_wire, --  input.wire
			output => cast207_output_wire        -- output.wire
		);

	cast208 : component alt_dspbuilder_cast_GNSB3OXIQS
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => memory_delay8_output_wire, --  input.wire
			output => cast208_output_wire        -- output.wire
		);

	cast209 : component alt_dspbuilder_cast_GN46N4UJ5S
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => comparator_result_wire, --  input.wire
			output => cast209_output_wire     -- output.wire
		);

	cast210 : component alt_dspbuilder_cast_GNXDXNUGW4
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => pixel_in_0_output_wire, --  input.wire
			output => cast210_output_wire     -- output.wire
		);

	cast211 : component alt_dspbuilder_cast_GN46N4UJ5S
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => comparator1_result_wire, --  input.wire
			output => cast211_output_wire      -- output.wire
		);

	cast212 : component alt_dspbuilder_cast_GN5D52DF5S
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => counter2_q_wire,     --  input.wire
			output => cast212_output_wire  -- output.wire
		);

	cast213 : component alt_dspbuilder_cast_GN46N4UJ5S
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => comparator3_result_wire, --  input.wire
			output => cast213_output_wire      -- output.wire
		);

	cast214 : component alt_dspbuilder_cast_GNRXYRYI2J
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => constant8_output_wire, --  input.wire
			output => cast214_output_wire    -- output.wire
		);

	cast215 : component alt_dspbuilder_cast_GNBKDIMZSI
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => constant9_output_wire, --  input.wire
			output => cast215_output_wire    -- output.wire
		);

	cast216 : component alt_dspbuilder_cast_GN46N4UJ5S
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => comparator7_result_wire, --  input.wire
			output => cast216_output_wire      -- output.wire
		);

	cast217 : component alt_dspbuilder_cast_GN46N4UJ5S
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => comparator7_result_wire, --  input.wire
			output => cast217_output_wire      -- output.wire
		);

	cast218 : component alt_dspbuilder_cast_GNNDZ2WJEB
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => memory_delay1_output_wire, --  input.wire
			output => cast218_output_wire        -- output.wire
		);

	cast219 : component alt_dspbuilder_cast_GN46N4UJ5S
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => comparator7_result_wire, --  input.wire
			output => cast219_output_wire      -- output.wire
		);

	cast220 : component alt_dspbuilder_cast_GNOZDXZSET
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => multiplexer4_result_wire, --  input.wire
			output => cast220_output_wire       -- output.wire
		);

	cast221 : component alt_dspbuilder_cast_GNACWQQVMS
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => histogram_q_wire,    --  input.wire
			output => cast221_output_wire  -- output.wire
		);

	cast222 : component alt_dspbuilder_cast_GNOZDXZSET
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => memory_delay5_output_wire, --  input.wire
			output => cast222_output_wire        -- output.wire
		);

	cast223 : component alt_dspbuilder_cast_GNQ4YFQS5C
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => histogram_q_wire,    --  input.wire
			output => cast223_output_wire  -- output.wire
		);

	cast224 : component alt_dspbuilder_cast_GNJYJUBV3U
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => multiplexer2_result_wire, --  input.wire
			output => cast224_output_wire       -- output.wire
		);

	cast225 : component alt_dspbuilder_cast_GN5PMHXBFJ
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => multiplexer7_result_wire, --  input.wire
			output => cast225_output_wire       -- output.wire
		);

	cast226 : component alt_dspbuilder_cast_GNZEACPTPO
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => multiplier1_result_wire, --  input.wire
			output => cast226_output_wire      -- output.wire
		);

	cast227 : component alt_dspbuilder_cast_GNNQZKMK3E
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => multiplexer3_result_wire, --  input.wire
			output => cast227_output_wire       -- output.wire
		);

	cast228 : component alt_dspbuilder_cast_GN5UGBMOKS
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => pipelined_adder1_result_wire, --  input.wire
			output => cast228_output_wire           -- output.wire
		);

	cast229 : component alt_dspbuilder_cast_GNSR6E4BZE
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => pipelined_adder1_result_wire, --  input.wire
			output => cast229_output_wire           -- output.wire
		);

	cast230 : component alt_dspbuilder_cast_GNDTOV7QCB
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => multiplexer2_result_wire, --  input.wire
			output => cast230_output_wire       -- output.wire
		);

	cast231 : component alt_dspbuilder_cast_GNAMS3PPNH
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => pipelined_adder2_result_wire, --  input.wire
			output => cast231_output_wire           -- output.wire
		);

	cast232 : component alt_dspbuilder_cast_GN46N4UJ5S
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => vcc_output_wire,     --  input.wire
			output => cast232_output_wire  -- output.wire
		);

end architecture rtl; -- of localedgepreserve_GN_localedgepreserve_Fusion_Cal_Weight
