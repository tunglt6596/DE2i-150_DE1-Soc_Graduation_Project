-- localedgepreserve_GN.vhd

-- Generated using ACDS version 17.1 590

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity localedgepreserve_GN is
	port (
		sink1_valid  : in  std_logic                    := '0';             --  sink1_valid.wire
		sink2_eop    : in  std_logic                    := '0';             --    sink2_eop.wire
		source_ready : in  std_logic                    := '0';             -- source_ready.wire
		source_data  : out std_logic_vector(7 downto 0);                    --  source_data.wire
		sink1_eop    : in  std_logic                    := '0';             --    sink1_eop.wire
		sink1_ready  : out std_logic;                                       --  sink1_ready.wire
		sink2_data   : in  std_logic_vector(7 downto 0) := (others => '0'); --   sink2_data.wire
		sink2_valid  : in  std_logic                    := '0';             --  sink2_valid.wire
		sink1_data   : in  std_logic_vector(7 downto 0) := (others => '0'); --   sink1_data.wire
		Clock        : in  std_logic                    := '0';             --        Clock.clk
		reset        : in  std_logic                    := '0';             --             .reset
		source_eop   : out std_logic;                                       --   source_eop.wire
		source_valid : out std_logic;                                       -- source_valid.wire
		source_sop   : out std_logic;                                       --   source_sop.wire
		sink2_sop    : in  std_logic                    := '0';             --    sink2_sop.wire
		sink1_sop    : in  std_logic                    := '0';             --    sink1_sop.wire
		sink2_ready  : out std_logic                                        --  sink2_ready.wire
	);
end entity localedgepreserve_GN;

architecture rtl of localedgepreserve_GN is
	component alt_dspbuilder_clock_GNN7TLRCSZ is
		port (
			aclr      : in  std_logic := 'X'; -- reset
			aclr_n    : in  std_logic := 'X'; -- reset_n
			aclr_out  : out std_logic;        -- reset
			clock     : in  std_logic := 'X'; -- clk
			clock_out : out std_logic         -- clk
		);
	end component alt_dspbuilder_clock_GNN7TLRCSZ;

	component alt_dspbuilder_port_GN37ALZBS4 is
		port (
			input  : in  std_logic := 'X'; -- wire
			output : out std_logic         -- wire
		);
	end component alt_dspbuilder_port_GN37ALZBS4;

	component alt_dspbuilder_multiplexer_GNIM5IEXF4 is
		generic (
			number_inputs          : natural  := 4;
			pipeline               : natural  := 0;
			width                  : positive := 8;
			HDLTYPE                : string   := "STD_LOGIC_VECTOR";
			use_one_hot_select_bus : natural  := 0
		);
		port (
			clock     : in  std_logic                    := 'X';             -- clk
			aclr      : in  std_logic                    := 'X';             -- reset
			sel       : in  std_logic_vector(0 downto 0) := (others => 'X'); -- wire
			result    : out std_logic_vector(8 downto 0);                    -- wire
			ena       : in  std_logic                    := 'X';             -- wire
			user_aclr : in  std_logic                    := 'X';             -- wire
			in0       : in  std_logic_vector(8 downto 0) := (others => 'X'); -- wire
			in1       : in  std_logic_vector(8 downto 0) := (others => 'X')  -- wire
		);
	end component alt_dspbuilder_multiplexer_GNIM5IEXF4;

	component alt_dspbuilder_gnd_GN is
		port (
			output : out std_logic   -- wire
		);
	end component alt_dspbuilder_gnd_GN;

	component alt_dspbuilder_vcc_GN is
		port (
			output : out std_logic   -- wire
		);
	end component alt_dspbuilder_vcc_GN;

	component alt_dspbuilder_comparator_GN is
		generic (
			Operator  : string  := "Altaeb";
			lpm_width : natural := 8
		);
		port (
			clock  : in  std_logic                              := 'X';             -- clk
			dataa  : in  std_logic_vector(lpm_width-1 downto 0) := (others => 'X'); -- wire
			datab  : in  std_logic_vector(lpm_width-1 downto 0) := (others => 'X'); -- wire
			result : out std_logic;                                                 -- wire
			sclr   : in  std_logic                              := 'X'              -- clk
		);
	end component alt_dspbuilder_comparator_GN;

	component alt_dspbuilder_extract_bit_GNN5FDHW3U is
		generic (
			ExtractedBit : natural := 0;
			width        : natural := 4
		);
		port (
			aclr   : in  std_logic                          := 'X';             -- clk
			clock  : in  std_logic                          := 'X';             -- clk
			input  : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			output : out std_logic                                              -- wire
		);
	end component alt_dspbuilder_extract_bit_GNN5FDHW3U;

	component localedgepreserve_GN_localedgepreserve_Fusion is
		port (
			pixel_out : out std_logic_vector(8 downto 0);                    -- wire
			pixel1_in : in  std_logic_vector(7 downto 0) := (others => 'X'); -- wire
			Clock     : in  std_logic                    := 'X';             -- clk
			reset     : in  std_logic                    := 'X';             -- reset
			valid2_in : in  std_logic                    := 'X';             -- wire
			sof_out   : out std_logic;                                       -- wire
			valid_out : out std_logic;                                       -- wire
			valid1_in : in  std_logic                    := 'X';             -- wire
			pixel2_in : in  std_logic_vector(7 downto 0) := (others => 'X'); -- wire
			eof_out   : out std_logic;                                       -- wire
			eof1_in   : in  std_logic                    := 'X';             -- wire
			eof2_in   : in  std_logic                    := 'X'              -- wire
		);
	end component localedgepreserve_GN_localedgepreserve_Fusion;

	component alt_dspbuilder_cast_GNMBFHMJNM is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(8 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(7 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNMBFHMJNM;

	component alt_dspbuilder_port_GNA5S4SQDN is
		port (
			input  : in  std_logic_vector(7 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(7 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNA5S4SQDN;

	component alt_dspbuilder_logical_bit_op_GNA5ZFEL7V is
		generic (
			LogicalOp     : string   := "AltAND";
			number_inputs : positive := 2
		);
		port (
			result : out std_logic;        -- wire
			data0  : in  std_logic := 'X'; -- wire
			data1  : in  std_logic := 'X'  -- wire
		);
	end component alt_dspbuilder_logical_bit_op_GNA5ZFEL7V;

	component alt_dspbuilder_constant_GNA4WR7CCY is
		generic (
			BitPattern : string  := "0000";
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(10 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GNA4WR7CCY;

	component alt_dspbuilder_constant_GNRT4BCWLZ is
		generic (
			BitPattern : string  := "0000";
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(8 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GNRT4BCWLZ;

	component alt_dspbuilder_bus_concat_GNMCLODSEX is
		generic (
			widthA : natural := 8;
			widthB : natural := 8
		);
		port (
			a      : in  std_logic_vector(widthA-1 downto 0)        := (others => 'X'); -- wire
			aclr   : in  std_logic                                  := 'X';             -- clk
			b      : in  std_logic_vector(widthB-1 downto 0)        := (others => 'X'); -- wire
			clock  : in  std_logic                                  := 'X';             -- clk
			output : out std_logic_vector(widthA+widthB-1 downto 0)                     -- wire
		);
	end component alt_dspbuilder_bus_concat_GNMCLODSEX;

	component alt_dspbuilder_fifo_GNC2APWQ5P is
		generic (
			numwords       : positive := 64;
			use_eab        : natural  := 1;
			ram_block_type : string   := "AUTO";
			width          : positive := 8;
			showahead_mode : natural  := 0;
			family         : string   := "Stratix"
		);
		port (
			clock : in  std_logic                     := 'X';             -- clk
			aclr  : in  std_logic                     := 'X';             -- reset
			data  : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- wire
			wrreq : in  std_logic                     := 'X';             -- wire
			rdreq : in  std_logic                     := 'X';             -- wire
			full  : out std_logic;                                        -- wire
			empty : out std_logic;                                        -- wire
			q     : out std_logic_vector(8 downto 0);                     -- wire
			usedw : out std_logic_vector(10 downto 0);                    -- wire
			sclr  : in  std_logic                     := 'X'              -- wire
		);
	end component alt_dspbuilder_fifo_GNC2APWQ5P;

	component alt_dspbuilder_cast_GNZZO4R4AV is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(10 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(11 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNZZO4R4AV;

	component alt_dspbuilder_cast_GN46N4UJ5S is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic                    := 'X'; -- wire
			output : out std_logic_vector(0 downto 0)         -- wire
		);
	end component alt_dspbuilder_cast_GN46N4UJ5S;

	signal multiplexeruser_aclrgnd_output_wire       : std_logic;                     -- Multiplexeruser_aclrGND:output -> Multiplexer:user_aclr
	signal multiplexerenavcc_output_wire             : std_logic;                     -- MultiplexerenaVCC:output -> Multiplexer:ena
	signal multiplexer1user_aclrgnd_output_wire      : std_logic;                     -- Multiplexer1user_aclrGND:output -> Multiplexer1:user_aclr
	signal multiplexer1enavcc_output_wire            : std_logic;                     -- Multiplexer1enaVCC:output -> Multiplexer1:ena
	signal fifo_1sclrgnd_output_wire                 : std_logic;                     -- FIFO_1sclrGND:output -> FIFO_1:sclr
	signal fifo_2sclrgnd_output_wire                 : std_logic;                     -- FIFO_2sclrGND:output -> FIFO_2:sclr
	signal bus_concatenation_output_wire             : std_logic_vector(8 downto 0);  -- Bus_Concatenation:output -> FIFO_1:data
	signal bus_concatenation1_output_wire            : std_logic_vector(8 downto 0);  -- Bus_Concatenation1:output -> FIFO_2:data
	signal logical_bit_operator1_result_wire         : std_logic;                     -- Logical_Bit_Operator1:result -> [FIFO_1:rdreq, FIFO_2:rdreq, cast324:input, cast325:input, localedgepreserve_Fusion_0:valid1_in, localedgepreserve_Fusion_0:valid2_in]
	signal bus_conversion_output_wire                : std_logic_vector(7 downto 0);  -- Bus_Conversion:output -> localedgepreserve_Fusion_0:pixel1_in
	signal extract_bit_output_wire                   : std_logic;                     -- Extract_Bit:output -> localedgepreserve_Fusion_0:eof1_in
	signal bus_conversion1_output_wire               : std_logic_vector(7 downto 0);  -- Bus_Conversion1:output -> localedgepreserve_Fusion_0:pixel2_in
	signal extract_bit1_output_wire                  : std_logic;                     -- Extract_Bit1:output -> localedgepreserve_Fusion_0:eof2_in
	signal comparator_result_wire                    : std_logic;                     -- Comparator:result -> Logical_Bit_Operator1:data0
	signal comparator1_result_wire                   : std_logic;                     -- Comparator1:result -> Logical_Bit_Operator1:data1
	signal constant_1_output_wire                    : std_logic_vector(8 downto 0);  -- Constant_1:output -> Multiplexer:in0
	signal fifo_1_q_wire                             : std_logic_vector(8 downto 0);  -- FIFO_1:q -> Multiplexer:in1
	signal multiplexer_result_wire                   : std_logic_vector(8 downto 0);  -- Multiplexer:result -> [Bus_Conversion:input, Extract_Bit:input]
	signal constant1_output_wire                     : std_logic_vector(8 downto 0);  -- Constant1:output -> Multiplexer1:in0
	signal fifo_2_q_wire                             : std_logic_vector(8 downto 0);  -- FIFO_2:q -> Multiplexer1:in1
	signal multiplexer1_result_wire                  : std_logic_vector(8 downto 0);  -- Multiplexer1:result -> [Bus_Conversion1:input, Extract_Bit1:input]
	signal sink1_data_0_output_wire                  : std_logic_vector(7 downto 0);  -- sink1_data_0:output -> Bus_Concatenation:b
	signal vcc3_output_wire                          : std_logic;                     -- VCC3:output -> sink1_ready_0:input
	signal sink1_valid_0_output_wire                 : std_logic;                     -- sink1_valid_0:output -> FIFO_1:wrreq
	signal sink2_data_0_output_wire                  : std_logic_vector(7 downto 0);  -- sink2_data_0:output -> Bus_Concatenation1:b
	signal vcc1_output_wire                          : std_logic;                     -- VCC1:output -> sink2_ready_0:input
	signal sink2_valid_0_output_wire                 : std_logic;                     -- sink2_valid_0:output -> FIFO_2:wrreq
	signal localedgepreserve_fusion_0_eof_out_wire   : std_logic;                     -- localedgepreserve_Fusion_0:eof_out -> source_eop_0:input
	signal localedgepreserve_fusion_0_sof_out_wire   : std_logic;                     -- localedgepreserve_Fusion_0:sof_out -> source_sop_0:input
	signal localedgepreserve_fusion_0_valid_out_wire : std_logic;                     -- localedgepreserve_Fusion_0:valid_out -> source_valid_0:input
	signal constant2_output_wire                     : std_logic_vector(10 downto 0); -- Constant2:output -> cast320:input
	signal cast320_output_wire                       : std_logic_vector(11 downto 0); -- cast320:output -> Comparator:datab
	signal constant3_output_wire                     : std_logic_vector(10 downto 0); -- Constant3:output -> cast321:input
	signal cast321_output_wire                       : std_logic_vector(11 downto 0); -- cast321:output -> Comparator1:datab
	signal fifo_1_usedw_wire                         : std_logic_vector(10 downto 0); -- FIFO_1:usedw -> cast322:input
	signal cast322_output_wire                       : std_logic_vector(11 downto 0); -- cast322:output -> Comparator:dataa
	signal fifo_2_usedw_wire                         : std_logic_vector(10 downto 0); -- FIFO_2:usedw -> cast323:input
	signal cast323_output_wire                       : std_logic_vector(11 downto 0); -- cast323:output -> Comparator1:dataa
	signal cast324_output_wire                       : std_logic_vector(0 downto 0);  -- cast324:output -> Multiplexer:sel
	signal cast325_output_wire                       : std_logic_vector(0 downto 0);  -- cast325:output -> Multiplexer1:sel
	signal sink1_eop_0_output_wire                   : std_logic;                     -- sink1_eop_0:output -> cast326:input
	signal cast326_output_wire                       : std_logic_vector(0 downto 0);  -- cast326:output -> Bus_Concatenation:a
	signal sink2_eop_0_output_wire                   : std_logic;                     -- sink2_eop_0:output -> cast327:input
	signal cast327_output_wire                       : std_logic_vector(0 downto 0);  -- cast327:output -> Bus_Concatenation1:a
	signal localedgepreserve_fusion_0_pixel_out_wire : std_logic_vector(8 downto 0);  -- localedgepreserve_Fusion_0:pixel_out -> cast328:input
	signal cast328_output_wire                       : std_logic_vector(7 downto 0);  -- cast328:output -> source_data_0:input
	signal clock_0_clock_output_clk                  : std_logic;                     -- Clock_0:clock_out -> [Bus_Concatenation1:clock, Bus_Concatenation:clock, Comparator1:clock, Comparator:clock, Extract_Bit1:clock, Extract_Bit:clock, FIFO_1:clock, FIFO_2:clock, Multiplexer1:clock, Multiplexer:clock, localedgepreserve_Fusion_0:Clock]
	signal clock_0_clock_output_reset                : std_logic;                     -- Clock_0:aclr_out -> [Bus_Concatenation1:aclr, Bus_Concatenation:aclr, Comparator1:sclr, Comparator:sclr, Extract_Bit1:aclr, Extract_Bit:aclr, FIFO_1:aclr, FIFO_2:aclr, Multiplexer1:aclr, Multiplexer:aclr, localedgepreserve_Fusion_0:reset]

begin

	clock_0 : component alt_dspbuilder_clock_GNN7TLRCSZ
		port map (
			clock_out => clock_0_clock_output_clk,   -- clock_output.clk
			aclr_out  => clock_0_clock_output_reset, --             .reset
			clock     => Clock,                      --        clock.clk
			aclr      => reset                       --             .reset
		);

	source_ready_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => source_ready, --  input.wire
			output => open          -- output.wire
		);

	multiplexer : component alt_dspbuilder_multiplexer_GNIM5IEXF4
		generic map (
			number_inputs          => 2,
			pipeline               => 0,
			width                  => 9,
			HDLTYPE                => "STD_LOGIC_VECTOR",
			use_one_hot_select_bus => 0
		)
		port map (
			clock     => clock_0_clock_output_clk,            -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,          --           .reset
			sel       => cast324_output_wire,                 --        sel.wire
			result    => multiplexer_result_wire,             --     result.wire
			ena       => multiplexerenavcc_output_wire,       --        ena.wire
			user_aclr => multiplexeruser_aclrgnd_output_wire, --  user_aclr.wire
			in0       => constant_1_output_wire,              --        in0.wire
			in1       => fifo_1_q_wire                        --        in1.wire
		);

	multiplexeruser_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplexeruser_aclrgnd_output_wire  -- output.wire
		);

	multiplexerenavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => multiplexerenavcc_output_wire  -- output.wire
		);

	sink2_ready_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => vcc1_output_wire, --  input.wire
			output => sink2_ready       -- output.wire
		);

	comparator : component alt_dspbuilder_comparator_GN
		generic map (
			Operator  => "Altagb",
			lpm_width => 12
		)
		port map (
			clock  => clock_0_clock_output_clk,   -- clock_sclr.clk
			sclr   => clock_0_clock_output_reset, --           .reset
			dataa  => cast322_output_wire,        --      dataa.wire
			datab  => cast320_output_wire,        --      datab.wire
			result => comparator_result_wire      --     result.wire
		);

	vcc1 : component alt_dspbuilder_vcc_GN
		port map (
			output => vcc1_output_wire  -- output.wire
		);

	vcc3 : component alt_dspbuilder_vcc_GN
		port map (
			output => vcc3_output_wire  -- output.wire
		);

	extract_bit : component alt_dspbuilder_extract_bit_GNN5FDHW3U
		generic map (
			ExtractedBit => 8,
			width        => 9
		)
		port map (
			clock  => clock_0_clock_output_clk,   -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset, --           .reset
			input  => multiplexer_result_wire,    --      input.wire
			output => extract_bit_output_wire     --     output.wire
		);

	sink2_valid_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => sink2_valid,               --  input.wire
			output => sink2_valid_0_output_wire  -- output.wire
		);

	localedgepreserve_fusion_0 : component localedgepreserve_GN_localedgepreserve_Fusion
		port map (
			pixel_out => localedgepreserve_fusion_0_pixel_out_wire, -- pixel_out.wire
			pixel1_in => bus_conversion_output_wire,                -- pixel1_in.wire
			Clock     => clock_0_clock_output_clk,                  --     Clock.clk
			reset     => clock_0_clock_output_reset,                --          .reset
			valid2_in => logical_bit_operator1_result_wire,         -- valid2_in.wire
			sof_out   => localedgepreserve_fusion_0_sof_out_wire,   --   sof_out.wire
			valid_out => localedgepreserve_fusion_0_valid_out_wire, -- valid_out.wire
			valid1_in => logical_bit_operator1_result_wire,         -- valid1_in.wire
			pixel2_in => bus_conversion1_output_wire,               -- pixel2_in.wire
			eof_out   => localedgepreserve_fusion_0_eof_out_wire,   --   eof_out.wire
			eof1_in   => extract_bit_output_wire,                   --   eof1_in.wire
			eof2_in   => extract_bit1_output_wire                   --   eof2_in.wire
		);

	bus_conversion : component alt_dspbuilder_cast_GNMBFHMJNM
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => multiplexer_result_wire,    --  input.wire
			output => bus_conversion_output_wire  -- output.wire
		);

	bus_conversion1 : component alt_dspbuilder_cast_GNMBFHMJNM
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => multiplexer1_result_wire,    --  input.wire
			output => bus_conversion1_output_wire  -- output.wire
		);

	source_data_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => cast328_output_wire, --  input.wire
			output => source_data          -- output.wire
		);

	logical_bit_operator1 : component alt_dspbuilder_logical_bit_op_GNA5ZFEL7V
		generic map (
			LogicalOp     => "AltAND",
			number_inputs => 2
		)
		port map (
			result => logical_bit_operator1_result_wire, -- result.wire
			data0  => comparator_result_wire,            --  data0.wire
			data1  => comparator1_result_wire            --  data1.wire
		);

	sink1_ready_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => vcc3_output_wire, --  input.wire
			output => sink1_ready       -- output.wire
		);

	source_eop_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => localedgepreserve_fusion_0_eof_out_wire, --  input.wire
			output => source_eop                               -- output.wire
		);

	constant2 : component alt_dspbuilder_constant_GNA4WR7CCY
		generic map (
			BitPattern => "00001100011",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 11
		)
		port map (
			output => constant2_output_wire  -- output.wire
		);

	constant3 : component alt_dspbuilder_constant_GNA4WR7CCY
		generic map (
			BitPattern => "00001100011",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 11
		)
		port map (
			output => constant3_output_wire  -- output.wire
		);

	constant1 : component alt_dspbuilder_constant_GNRT4BCWLZ
		generic map (
			BitPattern => "000000000",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 9
		)
		port map (
			output => constant1_output_wire  -- output.wire
		);

	sink2_data_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => sink2_data,               --  input.wire
			output => sink2_data_0_output_wire  -- output.wire
		);

	sink1_sop_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => sink1_sop, --  input.wire
			output => open       -- output.wire
		);

	bus_concatenation1 : component alt_dspbuilder_bus_concat_GNMCLODSEX
		generic map (
			widthA => 1,
			widthB => 8
		)
		port map (
			clock  => clock_0_clock_output_clk,       -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,     --           .reset
			a      => cast327_output_wire,            --          a.wire
			b      => sink2_data_0_output_wire,       --          b.wire
			output => bus_concatenation1_output_wire  --     output.wire
		);

	source_sop_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => localedgepreserve_fusion_0_sof_out_wire, --  input.wire
			output => source_sop                               -- output.wire
		);

	sink1_eop_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => sink1_eop,               --  input.wire
			output => sink1_eop_0_output_wire  -- output.wire
		);

	sink1_valid_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => sink1_valid,               --  input.wire
			output => sink1_valid_0_output_wire  -- output.wire
		);

	bus_concatenation : component alt_dspbuilder_bus_concat_GNMCLODSEX
		generic map (
			widthA => 1,
			widthB => 8
		)
		port map (
			clock  => clock_0_clock_output_clk,      -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,    --           .reset
			a      => cast326_output_wire,           --          a.wire
			b      => sink1_data_0_output_wire,      --          b.wire
			output => bus_concatenation_output_wire  --     output.wire
		);

	multiplexer1 : component alt_dspbuilder_multiplexer_GNIM5IEXF4
		generic map (
			number_inputs          => 2,
			pipeline               => 0,
			width                  => 9,
			HDLTYPE                => "STD_LOGIC_VECTOR",
			use_one_hot_select_bus => 0
		)
		port map (
			clock     => clock_0_clock_output_clk,             -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,           --           .reset
			sel       => cast325_output_wire,                  --        sel.wire
			result    => multiplexer1_result_wire,             --     result.wire
			ena       => multiplexer1enavcc_output_wire,       --        ena.wire
			user_aclr => multiplexer1user_aclrgnd_output_wire, --  user_aclr.wire
			in0       => constant1_output_wire,                --        in0.wire
			in1       => fifo_2_q_wire                         --        in1.wire
		);

	multiplexer1user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplexer1user_aclrgnd_output_wire  -- output.wire
		);

	multiplexer1enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => multiplexer1enavcc_output_wire  -- output.wire
		);

	sink2_eop_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => sink2_eop,               --  input.wire
			output => sink2_eop_0_output_wire  -- output.wire
		);

	comparator1 : component alt_dspbuilder_comparator_GN
		generic map (
			Operator  => "Altagb",
			lpm_width => 12
		)
		port map (
			clock  => clock_0_clock_output_clk,   -- clock_sclr.clk
			sclr   => clock_0_clock_output_reset, --           .reset
			dataa  => cast323_output_wire,        --      dataa.wire
			datab  => cast321_output_wire,        --      datab.wire
			result => comparator1_result_wire     --     result.wire
		);

	sink1_data_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => sink1_data,               --  input.wire
			output => sink1_data_0_output_wire  -- output.wire
		);

	sink2_sop_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => sink2_sop, --  input.wire
			output => open       -- output.wire
		);

	fifo_1 : component alt_dspbuilder_fifo_GNC2APWQ5P
		generic map (
			numwords       => 2048,
			use_eab        => 1,
			ram_block_type => "AUTO",
			width          => 9,
			showahead_mode => 0,
			family         => "Cyclone V"
		)
		port map (
			clock => clock_0_clock_output_clk,          -- clock_aclr.clk
			aclr  => clock_0_clock_output_reset,        --           .reset
			data  => bus_concatenation_output_wire,     --       data.wire
			wrreq => sink1_valid_0_output_wire,         --      wrreq.wire
			rdreq => logical_bit_operator1_result_wire, --      rdreq.wire
			full  => open,                              --       full.wire
			empty => open,                              --      empty.wire
			q     => fifo_1_q_wire,                     --          q.wire
			usedw => fifo_1_usedw_wire,                 --      usedw.wire
			sclr  => fifo_1sclrgnd_output_wire          --       sclr.wire
		);

	fifo_1sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => fifo_1sclrgnd_output_wire  -- output.wire
		);

	fifo_2 : component alt_dspbuilder_fifo_GNC2APWQ5P
		generic map (
			numwords       => 2048,
			use_eab        => 1,
			ram_block_type => "AUTO",
			width          => 9,
			showahead_mode => 0,
			family         => "Cyclone V"
		)
		port map (
			clock => clock_0_clock_output_clk,          -- clock_aclr.clk
			aclr  => clock_0_clock_output_reset,        --           .reset
			data  => bus_concatenation1_output_wire,    --       data.wire
			wrreq => sink2_valid_0_output_wire,         --      wrreq.wire
			rdreq => logical_bit_operator1_result_wire, --      rdreq.wire
			full  => open,                              --       full.wire
			empty => open,                              --      empty.wire
			q     => fifo_2_q_wire,                     --          q.wire
			usedw => fifo_2_usedw_wire,                 --      usedw.wire
			sclr  => fifo_2sclrgnd_output_wire          --       sclr.wire
		);

	fifo_2sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => fifo_2sclrgnd_output_wire  -- output.wire
		);

	source_valid_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => localedgepreserve_fusion_0_valid_out_wire, --  input.wire
			output => source_valid                               -- output.wire
		);

	constant_1 : component alt_dspbuilder_constant_GNRT4BCWLZ
		generic map (
			BitPattern => "000000000",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 9
		)
		port map (
			output => constant_1_output_wire  -- output.wire
		);

	extract_bit1 : component alt_dspbuilder_extract_bit_GNN5FDHW3U
		generic map (
			ExtractedBit => 8,
			width        => 9
		)
		port map (
			clock  => clock_0_clock_output_clk,   -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset, --           .reset
			input  => multiplexer1_result_wire,   --      input.wire
			output => extract_bit1_output_wire    --     output.wire
		);

	cast320 : component alt_dspbuilder_cast_GNZZO4R4AV
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => constant2_output_wire, --  input.wire
			output => cast320_output_wire    -- output.wire
		);

	cast321 : component alt_dspbuilder_cast_GNZZO4R4AV
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => constant3_output_wire, --  input.wire
			output => cast321_output_wire    -- output.wire
		);

	cast322 : component alt_dspbuilder_cast_GNZZO4R4AV
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => fifo_1_usedw_wire,   --  input.wire
			output => cast322_output_wire  -- output.wire
		);

	cast323 : component alt_dspbuilder_cast_GNZZO4R4AV
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => fifo_2_usedw_wire,   --  input.wire
			output => cast323_output_wire  -- output.wire
		);

	cast324 : component alt_dspbuilder_cast_GN46N4UJ5S
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => logical_bit_operator1_result_wire, --  input.wire
			output => cast324_output_wire                -- output.wire
		);

	cast325 : component alt_dspbuilder_cast_GN46N4UJ5S
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => logical_bit_operator1_result_wire, --  input.wire
			output => cast325_output_wire                -- output.wire
		);

	cast326 : component alt_dspbuilder_cast_GN46N4UJ5S
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => sink1_eop_0_output_wire, --  input.wire
			output => cast326_output_wire      -- output.wire
		);

	cast327 : component alt_dspbuilder_cast_GN46N4UJ5S
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => sink2_eop_0_output_wire, --  input.wire
			output => cast327_output_wire      -- output.wire
		);

	cast328 : component alt_dspbuilder_cast_GNMBFHMJNM
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => localedgepreserve_fusion_0_pixel_out_wire, --  input.wire
			output => cast328_output_wire                        -- output.wire
		);

end architecture rtl; -- of localedgepreserve_GN
